module FNIRSI_1014D
(
  output wire io_i2c_scl,
  inout wire io_i2c_sda,
  input wire i_clk2,
  input wire i_clk1,
  output wire o_pwm_display,
  input wire i_mcu_rws,
  input wire i_mcu_dcs,
  input wire i_mcu_clk,
  output wire o_dac_d[1],
  output wire o_dac_d[0],
  inout wire io_mcu_d[4],
  inout wire io_mcu_d[5],
  inout wire io_mcu_d[6],
  inout wire io_mcu_d[7],
  output wire o_dac_d[2],
  output wire o_dac_d[5],
  output wire o_dac_d[3],
  output wire o_dac_d[4],
  inout wire io_mcu_d[2],
  inout wire io_mcu_d[3],
  inout wire io_mcu_d[1],
  inout wire io_mcu_d[0],
  output wire o_dac_d[6],
  output wire o_dac_d[7],
  output wire o_ac_dc_2,
  output wire o_ac_dc_1,
  output wire o_relay1_2,
  output wire o_relay1_1,
  output wire o_relay2_2,
  output wire o_relay1_3,
  output wire o_relay2_3,
  output wire o_relay2_1,
  input wire i_adc1B_d[6],
  output wire o_adc1_encB,
  input wire i_adc1B_d[7],
  input wire i_adc2A_d[6],
  input wire i_adc2A_d[5],
  output wire o_adc2_encA,
  input wire i_adc2A_d[7],
  input wire i_adc2A_d[3],
  input wire i_adc2A_d[4],
  input wire i_adc1B_d[2],
  input wire i_adc1B_d[3],
  input wire i_adc1B_d[4],
  input wire i_adc1B_d[5],
  input wire i_adc2A_d[0],
  input wire i_adc2A_d[1],
  input wire i_adc2A_d[2],
  input wire i_adc1B_d[0],
  input wire i_adc1B_d[1],
  input wire i_adc2B_d[1],
  input wire i_adc2B_d[0],
  input wire i_adc2B_d[2],
  input wire i_adc2B_d[4],
  input wire i_adc2B_d[3],
  input wire i_adc2B_d[5],
  input wire i_adc2B_d[6],
  output wire o_adc2_encB,
  input wire i_adc2B_d[7],
  output wire o_offset_2,
  output wire o_offset_1,
  output wire o_adc1_encA,
  input wire i_adc1A_d[7],
  input wire i_adc1A_d[5],
  input wire i_adc1A_d[6],
  input wire i_adc1A_d[3],
  input wire i_adc1A_d[4],
  input wire i_adc1A_d[2],
  input wire i_adc1A_d[0],
  input wire i_adc1A_d[1]
);

  assign io_i2c_scl = net_341;
  assign io_i2c_sda = net_194 ? net_342 : 1'bZ;
  assign o_pwm_display = net_1118;
  assign o_dac_d[1] = net_23;
  assign o_dac_d[0] = net_22;
  assign io_mcu_d[4] = net_288 ? net_324 : 1'bZ;
  assign io_mcu_d[5] = net_288 ? net_256 : 1'bZ;
  assign io_mcu_d[6] = net_288 ? net_190 : 1'bZ;
  assign io_mcu_d[7] = net_288 ? net_188 : 1'bZ;
  assign o_dac_d[2] = net_21;
  assign o_dac_d[5] = net_26;
  assign o_dac_d[3] = net_24;
  assign o_dac_d[4] = net_27;
  assign io_mcu_d[2] = net_288 ? net_908 : 1'bZ;
  assign io_mcu_d[3] = net_288 ? net_262 : 1'bZ;
  assign io_mcu_d[1] = net_288 ? net_662 : 1'bZ;
  assign io_mcu_d[0] = net_288 ? net_911 : 1'bZ;
  assign o_dac_d[6] = net_25;
  assign o_dac_d[7] = net_28;
  assign o_ac_dc_2 = net_253;
  assign o_ac_dc_1 = net_322;
  assign o_relay1_2 = net_866;
  assign o_relay1_1 = net_864;
  assign o_relay2_2 = net_972;
  assign o_relay1_3 = net_865;
  assign o_relay2_3 = net_973;
  assign o_relay2_1 = net_971;
  assign o_adc1_encB = net_1502;
  assign o_adc2_encA = net_1471;
  assign o_adc2_encB = net_1472;
  assign o_offset_2 = net_788;
  assign o_offset_1 = net_990;
  assign o_adc1_encA = net_1618;

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hEEAA"),
    .INIT_LUTG0("16'hCC00"),
    .INIT_LUTF1("16'h00AA"),
    .INIT_LUTG1("16'hCCEE"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_101
  (
    .clk(gclk_9),
    .a({net_66,net_65}),
    .b({net_512,net_121}),
    .d({net_234,net_512}),
    .e({net_123,net_234}),
    .q({net_66,net_65})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h000A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD_CARRY"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("F"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_102
  (
    .clk(gclk_7),
    .sr(net_137),
    .a({net_68,1'b0}),
    .q({net_68,open_n0}),
    .fco(block_102_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_103
  (
    .clk(gclk_7),
    .sr(net_137),
    .a({net_67,net_69}),
    .b({1'b0,1'b0}),
    .fci(block_102_carry),
    .q({net_67,net_69}),
    .fco(block_103_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_104
  (
    .clk(gclk_7),
    .sr(net_137),
    .a({net_71,net_73}),
    .b({1'b0,1'b0}),
    .fci(block_103_carry),
    .q({net_71,net_73}),
    .fco(block_104_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_105
  (
    .clk(gclk_7),
    .sr(net_137),
    .a({net_70,net_72}),
    .b({1'b0,1'b0}),
    .fci(block_104_carry),
    .q({net_70,net_72}),
    .fco(block_105_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_106
  (
    .clk(gclk_7),
    .sr(net_137),
    .a({net_74,net_77}),
    .b({1'b0,1'b0}),
    .fci(block_105_carry),
    .q({net_74,net_77}),
    .fco(block_106_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_108
  (
    .clk(gclk_7),
    .sr(net_137),
    .a({open_n1,net_76}),
    .b({open_n2,1'b0}),
    .fci(block_106_carry),
    .q({open_n3,net_76})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hCF8E"),
    .INIT_LUTG0("16'h8E0C"),
    .INIT_LUTF1("16'h2302"),
    .INIT_LUTG1("16'hBF3B"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_107
  (
    .clk(gclk_9),
    .ce(net_221),
    .a({net_75,net_78}),
    .b({net_72,net_226}),
    .c({net_71,net_77}),
    .d({net_133,net_80}),
    .e({net_227,net_70}),
    .mi({io_mcu_d[4],io_mcu_d[6]}),
    .f({net_78,net_79}),
    .q({net_75,net_80})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hBB0B"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'hFF55"),
    .INIT_LUTG1("16'hF050"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_109
  (
    .clk(gclk_9),
    .ce(net_235),
    .a({net_82,net_81}),
    .b({open_n4,net_155}),
    .c({net_176,net_239}),
    .d({net_239,net_82}),
    .e({net_141,net_148}),
    .mi({io_mcu_d[5],io_mcu_d[4]}),
    .f({net_83,net_84}),
    .q({net_82,net_81})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hAFCF"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_110
  (
    .a({net_46,net_46}),
    .b({net_37,net_37}),
    .c({net_189,net_189}),
    .d({net_1044,net_1044}),
    .mi({open_n5,net_187}),
    .fx({open_n6,net_85})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hAFCF"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_111
  (
    .a({net_39,net_39}),
    .b({net_31,net_31}),
    .c({net_1044,net_189}),
    .d({net_189,net_1044}),
    .mi({open_n7,net_93}),
    .fx({open_n8,net_86})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h00FF"),
    .INIT_LUTG0("16'h80FF"),
    .INIT_LUTF1("16'h0001"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_112
  (
    .clk(gclk_5),
    .sr(net_90),
    .a({net_87,net_165}),
    .b({net_162,net_233}),
    .c({net_166,net_178}),
    .d({net_88,net_89}),
    .e({net_174,net_240}),
    .mi({net_169,net_171}),
    .f({net_89,net_90}),
    .q({net_87,net_88})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h5F3F"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_113
  (
    .a({net_43,net_43}),
    .b({net_33,net_33}),
    .c({net_189,net_189}),
    .d({net_1044,net_1044}),
    .mi({open_n9,net_92}),
    .fx({open_n10,net_91})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hAFCF"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_114
  (
    .a({net_44,net_44}),
    .b({net_34,net_34}),
    .c({net_1044,net_189}),
    .d({net_189,net_1044}),
    .mi({open_n11,net_96}),
    .fx({open_n12,net_95})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h5151"),
    .INIT_LUTG0("16'h0101"),
    .INIT_LUTF1("16'h00AF"),
    .INIT_LUTG1("16'h0005"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_115
  (
    .a({net_1044,net_189}),
    .b({open_n13,net_48}),
    .c({net_54,net_1044}),
    .d({net_189,open_n14}),
    .e({net_62,net_57}),
    .f({net_96,net_94})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0A0C"),
    .INIT_LUTG0("16'h0A0C"),
    .INIT_LUTF1("16'h003F"),
    .INIT_LUTG1("16'h000C"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_116
  (
    .a({open_n15,net_58}),
    .b({net_1044,net_52}),
    .c({net_60,net_189}),
    .d({net_189,net_1044}),
    .e({net_49,open_n16}),
    .f({net_93,net_92})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h888A"),
    .INIT_LUTG0("16'h8F8A"),
    .INIT_LUTF1("16'h888A"),
    .INIT_LUTG1("16'h88FA"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_117
  (
    .clk(gclk_9),
    .a({net_97,net_98}),
    .b({net_793,net_793}),
    .c({net_264,i_mcu_dcs}),
    .d({i_mcu_dcs,net_264}),
    .e({io_mcu_d[3],io_mcu_d[2]}),
    .q({net_97,net_98})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hB0AA"),
    .INIT_LUTG0("16'hBBBB"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hAAAA"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_118
  (
    .clk(gclk_9),
    .a({net_648,net_99}),
    .b({open_n17,net_793}),
    .c({open_n18,io_mcu_d[5]}),
    .d({open_n19,net_100}),
    .e({i_mcu_rws,i_mcu_dcs}),
    .f({net_100,open_n20}),
    .q({open_n21,net_99})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hBBAA"),
    .INIT_LUTG0("16'hBBB0"),
    .INIT_LUTF1("16'h888A"),
    .INIT_LUTG1("16'h8F8A"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_119
  (
    .clk(gclk_9),
    .a({net_104,net_102}),
    .b({net_793,net_793}),
    .c({i_mcu_dcs,io_mcu_d[2]}),
    .d({net_816,i_mcu_dcs}),
    .e({io_mcu_d[3],net_816}),
    .q({net_104,net_102})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h888A"),
    .INIT_LUTG0("16'h8F8A"),
    .INIT_LUTF1("16'h888A"),
    .INIT_LUTG1("16'h8F8A"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_120
  (
    .clk(gclk_9),
    .a({net_101,net_103}),
    .b({net_793,net_793}),
    .c({i_mcu_dcs,i_mcu_dcs}),
    .d({net_816,net_816}),
    .e({io_mcu_d[4],io_mcu_d[5]}),
    .q({net_101,net_103})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h000A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD_CARRY"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_125
  (
    .clk(gclk_9),
    .a({net_115,1'b0}),
    .mi({open_n22,net_115}),
    .f({net_114,open_n23}),
    .q({open_n24,net_112}),
    .fco(block_125_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_127
  (
    .clk(gclk_9),
    .a({1'b0,net_290}),
    .b({net_216,1'b0}),
    .mi({net_216,net_290}),
    .fci(block_125_carry),
    .f({net_113,net_109}),
    .q({net_111,net_110}),
    .fco(block_127_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_128
  (
    .clk(gclk_9),
    .a({1'b0,1'b0}),
    .b({net_108,net_66}),
    .mi({net_108,net_66}),
    .fci(block_127_carry),
    .f({net_122,net_123}),
    .q({net_117,net_120}),
    .fco(block_128_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_130
  (
    .clk(gclk_9),
    .a({1'b0,1'b0}),
    .b({net_65,net_107}),
    .mi({net_65,net_107}),
    .fci(block_128_carry),
    .f({net_121,net_124}),
    .q({net_119,net_118}),
    .fco(block_130_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_131
  (
    .clk(gclk_9),
    .a({1'b0,net_217}),
    .b({net_291,1'b0}),
    .mi({net_291,net_217}),
    .fci(block_130_carry),
    .f({net_125,net_127}),
    .q({net_128,net_130}),
    .fco(block_131_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_132
  (
    .clk(gclk_9),
    .a({open_n25,net_116}),
    .b({open_n26,1'b0}),
    .mi({open_n27,net_116}),
    .fci(block_131_carry),
    .f({open_n28,net_129}),
    .q({open_n29,net_126})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h2222"),
    .INIT_LUTG0("16'hFF22"),
    .INIT_LUTF1("16'hEEAA"),
    .INIT_LUTG1("16'hCC00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_126
  (
    .clk(gclk_9),
    .a({net_108,net_107}),
    .b({net_122,net_234}),
    .d({net_512,net_512}),
    .e({net_234,net_124}),
    .q({net_108,net_107})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0A0A"),
    .INIT_LUTG0("16'hFF0A"),
    .INIT_LUTF1("16'h0A0A"),
    .INIT_LUTG1("16'hFF0A"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_129
  (
    .clk(gclk_9),
    .a({net_115,net_116}),
    .c({net_234,net_234}),
    .d({net_512,net_512}),
    .e({net_114,net_129}),
    .q({net_115,net_116})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hF371"),
    .INIT_LUTG0("16'h7130"),
    .INIT_LUTF1("16'hF5F5"),
    .INIT_LUTG1("16'hD4D4"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_133
  (
    .clk(gclk_9),
    .ce(net_221),
    .a({net_131,net_132}),
    .b({net_68,net_73}),
    .c({net_69,net_223}),
    .d({open_n30,net_134}),
    .e({net_225,net_67}),
    .mi({io_mcu_d[1],io_mcu_d[2]}),
    .f({net_132,net_133}),
    .q({net_131,net_134})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h444D"),
    .INIT_LUTG0("16'h4DDD"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hC0C0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_134
  (
    .clk(gclk_9),
    .ce(net_138),
    .a({open_n31,net_135}),
    .b({net_1283,net_76}),
    .c({net_220,net_79}),
    .d({open_n32,net_136}),
    .e({net_452,net_74}),
    .mi({io_mcu_d[0],io_mcu_d[1]}),
    .f({net_138,net_137}),
    .q({net_136,net_135})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hAFCF"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_135
  (
    .a({net_38,net_38}),
    .b({net_29,net_29}),
    .c({net_1044,net_189}),
    .d({net_189,net_1044}),
    .mi({open_n33,net_94}),
    .fx({open_n34,net_146})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h5D04"),
    .INIT_LUTG0("16'hFF55"),
    .INIT_LUTF1("16'h5050"),
    .INIT_LUTG1("16'h5050"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_136
  (
    .clk(gclk_9),
    .ce(net_235),
    .a({net_141,net_139}),
    .b({open_n35,net_83}),
    .c({net_176,net_84}),
    .d({open_n36,net_165}),
    .e({open_n37,net_145}),
    .mi({io_mcu_d[6],io_mcu_d[7]}),
    .f({net_145,net_144}),
    .q({net_141,net_139})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hAF23"),
    .INIT_LUTG0("16'h0A02"),
    .INIT_LUTF1("16'h5151"),
    .INIT_LUTG1("16'h5100"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_137
  (
    .clk(gclk_9),
    .ce(net_235),
    .a({net_143,net_140}),
    .b({net_142,net_149}),
    .c({net_149,net_238}),
    .d({net_155,net_142}),
    .e({net_81,net_175}),
    .mi({io_mcu_d[3],io_mcu_d[2]}),
    .f({net_148,net_143}),
    .q({net_142,net_140})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hAFCF"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_138
  (
    .a({net_45,net_45}),
    .b({net_36,net_36}),
    .c({net_189,net_189}),
    .d({net_1044,net_1044}),
    .mi({open_n38,net_218}),
    .fx({open_n39,net_147})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hAFCF"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_139
  (
    .a({net_40,net_40}),
    .b({net_32,net_32}),
    .c({net_1044,net_189}),
    .d({net_189,net_1044}),
    .mi({open_n40,net_185}),
    .fx({open_n41,net_160})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h000A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_140
  (
    .clk(gclk_5),
    .sr(net_90),
    .a({net_150,1'b0}),
    .b({net_175,net_151}),
    .c({1'b0,1'b0}),
    .d({1'b0,open_n42}),
    .e({1'b0,open_n43}),
    .mi({net_154,net_159}),
    .f({net_154,open_n44}),
    .fx({net_152,net_159}),
    .q({net_150,net_151}),
    .fco(sig_140_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_141
  (
    .clk(gclk_5),
    .sr(net_90),
    .a({net_239,net_149}),
    .b({net_176,net_155}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_156,net_158}),
    .fci(sig_140_carry),
    .f({net_157,net_158}),
    .fx({net_153,net_156}),
    .q({net_155,net_149}),
    .fco(sig_141_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_143
  (
    .clk(gclk_5),
    .sr(net_90),
    .a({net_178,net_165}),
    .b({net_163,net_233}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_168,net_173}),
    .fci(sig_141_carry),
    .f({net_164,net_168}),
    .fx({net_173,net_170}),
    .q({net_165,net_163}),
    .fco(sig_143_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_144
  (
    .clk(gclk_5),
    .sr(net_90),
    .a({net_88,net_162}),
    .b({net_87,net_166}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_167,net_172}),
    .fci(sig_143_carry),
    .f({net_171,net_172}),
    .fx({net_169,net_167}),
    .q({net_166,net_162}),
    .fco(sig_144_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_145
  (
    .clk(gclk_5),
    .sr(net_90),
    .a({open_n45,net_174}),
    .c({1'b0,1'b0}),
    .d({open_n46,1'b0}),
    .mi({net_152,net_177}),
    .fci(sig_144_carry),
    .f({open_n47,net_177}),
    .q({net_175,net_174})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hAFCF"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_142
  (
    .a({net_41,net_41}),
    .b({net_30,net_30}),
    .c({net_189,net_189}),
    .d({net_1044,net_1044}),
    .mi({open_n48,net_192}),
    .fx({open_n49,net_161})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hAFCF"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_146
  (
    .a({net_42,net_42}),
    .b({net_35,net_35}),
    .c({net_189,net_189}),
    .d({net_1044,net_1044}),
    .mi({open_n50,net_259}),
    .fx({open_n51,net_179})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_147
  (
    .clk(gclk_5),
    .sr(net_90),
    .mi({net_153,net_164}),
    .q({net_176,net_178})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hAA00"),
    .INIT_LUTG0("16'hAA00"),
    .INIT_LUTF1("16'h5555"),
    .INIT_LUTG1("16'h5555"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_148
  (
    .clk(gclk_9),
    .ce(net_184),
    .a({net_248,i_mcu_rws}),
    .d({open_n52,i_mcu_dcs}),
    .mi({io_mcu_d[1],io_mcu_d[0]}),
    .f({net_182,net_184}),
    .q({net_181,net_180})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0A0C"),
    .INIT_LUT1("16'h0503"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_149
  (
    .a({net_59,net_730}),
    .b({net_50,net_739}),
    .c({net_189,net_189}),
    .d({net_1044,net_1044}),
    .f({net_185,net_183})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h2200"),
    .INIT_LUTG0("16'h2233"),
    .INIT_LUTF1("16'h0555"),
    .INIT_LUTG1("16'h0050"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_150
  (
    .a({net_189,net_734}),
    .b({open_n53,net_189}),
    .c({net_1044,open_n54}),
    .d({net_64,net_1044}),
    .e({net_53,net_740}),
    .f({net_187,net_186})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0053"),
    .INIT_LUT1("16'hACAC"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("F"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_151
  (
    .clk(gclk_3),
    .a({net_1197,net_56}),
    .b({net_1288,net_47}),
    .c({net_527,net_1044}),
    .d({open_n55,net_189}),
    .f({net_193,net_192}),
    .q({net_189,open_n56})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hCC55"),
    .INIT_LUTG0("16'hF0F0"),
    .INIT_LUTF1("16'hC0CC"),
    .INIT_LUTG1("16'hC0CC"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_152
  (
    .clk(gclk_9),
    .a({open_n57,net_191}),
    .b({net_468,net_531}),
    .c({net_310,net_190}),
    .d({net_190,i_mcu_dcs}),
    .e({open_n58,i_mcu_rws}),
    .f({net_191,open_n59}),
    .q({open_n60,net_190})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hCC0F"),
    .INIT_LUT1("16'hFF00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_153
  (
    .clk(gclk_9),
    .a({net_339,net_188}),
    .b({net_314,net_314}),
    .c({i_mcu_dcs,net_339}),
    .d({net_188,i_mcu_dcs}),
    .mi({open_n61,i_mcu_rws}),
    .q({open_n62,net_188})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0A00"),
    .INIT_LUT1("16'hFF0B"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_154
  (
    .clk(gclk_9),
    .a({io_mcu_d[6],io_mcu_d[6]}),
    .b({net_264,net_793}),
    .c({i_mcu_dcs,i_mcu_dcs}),
    .d({net_793,net_264}),
    .mi({open_n63,net_196}),
    .q({open_n64,net_196})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h888A"),
    .INIT_LUTG0("16'h8F8A"),
    .INIT_LUTF1("16'h5F5F"),
    .INIT_LUTG1("16'h005F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_155
  (
    .clk(gclk_9),
    .a({net_97,net_195}),
    .b({open_n65,net_793}),
    .c({net_952,i_mcu_dcs}),
    .d({net_195,net_264}),
    .e({net_962,io_mcu_d[4]}),
    .f({net_197,open_n66}),
    .q({open_n67,net_195})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hAAFA"),
    .INIT_LUT1("16'h3232"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("INV"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_156
  (
    .clk(gclk_8),
    .ce(net_248),
    .a({net_247,net_194}),
    .b({net_569,net_350}),
    .c({net_350,net_247}),
    .d({net_194,net_569}),
    .mi({open_n68,net_578}),
    .q({open_n69,net_194})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h888A"),
    .INIT_LUTG0("16'h8F8A"),
    .INIT_LUTF1("16'h5F5F"),
    .INIT_LUTG1("16'h005F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_157
  (
    .clk(gclk_9),
    .a({net_585,net_198}),
    .b({open_n70,net_793}),
    .c({net_98,i_mcu_dcs}),
    .d({net_198,net_264}),
    .e({net_843,io_mcu_d[0]}),
    .f({net_199,open_n71}),
    .q({open_n72,net_198})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0A00"),
    .INIT_LUT1("16'hAFAB"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_158
  (
    .clk(gclk_9),
    .a({net_793,io_mcu_d[7]}),
    .b({net_264,net_793}),
    .c({i_mcu_dcs,i_mcu_dcs}),
    .d({io_mcu_d[7],net_264}),
    .mi({open_n73,net_205}),
    .q({open_n74,net_205})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hBBAA"),
    .INIT_LUTG0("16'hBBB0"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hECA0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_159
  (
    .clk(gclk_9),
    .a({net_862,net_200}),
    .b({net_952,net_793}),
    .c({net_99,io_mcu_d[2]}),
    .d({net_200,i_mcu_dcs}),
    .e({net_943,net_100}),
    .f({net_203,open_n75}),
    .q({open_n76,net_200})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h888A"),
    .INIT_LUTG0("16'h8F8A"),
    .INIT_LUTF1("16'h77FF"),
    .INIT_LUTG1("16'h070F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_160
  (
    .clk(gclk_9),
    .a({net_951,net_201}),
    .b({net_862,net_793}),
    .c({net_840,i_mcu_dcs}),
    .d({net_201,net_265}),
    .e({net_103,io_mcu_d[1]}),
    .f({net_204,open_n77}),
    .q({open_n78,net_201})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0A00"),
    .INIT_LUT1("16'hCECF"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_161
  (
    .clk(gclk_9),
    .a({io_mcu_d[6],io_mcu_d[6]}),
    .b({net_793,net_793}),
    .c({i_mcu_dcs,i_mcu_dcs}),
    .d({net_816,net_816}),
    .mi({open_n79,net_202}),
    .q({open_n80,net_202})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0A00"),
    .INIT_LUT1("16'hCFCD"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_162
  (
    .clk(gclk_9),
    .a({net_816,io_mcu_d[7]}),
    .b({net_793,net_793}),
    .c({i_mcu_dcs,i_mcu_dcs}),
    .d({io_mcu_d[7],net_816}),
    .mi({open_n81,net_207}),
    .q({open_n82,net_207})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h888A"),
    .INIT_LUTG0("16'h8F8A"),
    .INIT_LUTF1("16'h3F3F"),
    .INIT_LUTG1("16'h003F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_163
  (
    .clk(gclk_9),
    .a({open_n83,net_206}),
    .b({net_843,net_793}),
    .c({net_102,i_mcu_dcs}),
    .d({net_206,net_816}),
    .e({net_950,io_mcu_d[1]}),
    .f({net_209,open_n84}),
    .q({open_n85,net_206})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0A00"),
    .INIT_LUT1("16'hCECF"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_164
  (
    .clk(gclk_9),
    .a({io_mcu_d[5],io_mcu_d[5]}),
    .b({net_793,net_793}),
    .c({i_mcu_dcs,i_mcu_dcs}),
    .d({net_286,net_286}),
    .mi({open_n86,net_208}),
    .q({open_n87,net_208})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h888A"),
    .INIT_LUTG0("16'h8F8A"),
    .INIT_LUTF1("16'h5F5F"),
    .INIT_LUTG1("16'h005F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_165
  (
    .clk(gclk_9),
    .a({net_208,net_210}),
    .b({open_n88,net_793}),
    .c({net_843,i_mcu_dcs}),
    .d({net_210,net_286}),
    .e({net_863,io_mcu_d[2]}),
    .f({net_211,open_n89}),
    .q({open_n90,net_210})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hBBAA"),
    .INIT_LUTG0("16'hBBB0"),
    .INIT_LUTF1("16'h33FF"),
    .INIT_LUTG1("16'h1155"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_166
  (
    .clk(gclk_9),
    .a({net_564,net_212}),
    .b({net_668,net_793}),
    .c({open_n91,io_mcu_d[1]}),
    .d({net_212,i_mcu_dcs}),
    .e({net_214,net_286}),
    .f({net_213,open_n92}),
    .q({open_n93,net_212})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hBBAA"),
    .INIT_LUTG0("16'hBBB0"),
    .INIT_LUTF1("16'hBBAA"),
    .INIT_LUTG1("16'hBBB0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_167
  (
    .clk(gclk_9),
    .a({net_215,net_214}),
    .b({net_793,net_793}),
    .c({io_mcu_d[4],io_mcu_d[3]}),
    .d({i_mcu_dcs,i_mcu_dcs}),
    .e({net_100,net_100}),
    .q({net_215,net_214})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hCE0A"),
    .INIT_LUT1("16'hCE0A"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_172
  (
    .clk(gclk_9),
    .a({net_216,net_217}),
    .b({net_113,net_127}),
    .c({net_234,net_234}),
    .d({net_512,net_512}),
    .q({net_216,net_217})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0503"),
    .INIT_LUT1("16'h0053"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_173
  (
    .a({net_63,net_700}),
    .b({net_55,net_692}),
    .c({net_1044,net_189}),
    .d({net_189,net_1044}),
    .f({net_218,net_219})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'hCCCC"),
    .INIT_LUTF1("16'hC0C0"),
    .INIT_LUTG1("16'hC0C0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_174
  (
    .clk(gclk_9),
    .ce(net_221),
    .b({net_452,net_309}),
    .c({net_315,open_n94}),
    .e({open_n95,net_452}),
    .mi({io_mcu_d[5],io_mcu_d[7]}),
    .f({net_222,net_224}),
    .q({net_227,net_226})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h8000"),
    .INIT_LUT1("16'h8800"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_175
  (
    .clk(gclk_9),
    .ce(net_221),
    .a({net_220,net_308}),
    .b({net_452,net_316}),
    .c({open_n96,net_180}),
    .d({net_1141,net_181}),
    .mi({io_mcu_d[0],io_mcu_d[3]}),
    .f({net_221,net_220}),
    .q({net_225,net_223})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h8800"),
    .INIT_LUT1("16'hD4DD"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_176
  (
    .clk(gclk_9),
    .ce(net_235),
    .a({net_229,net_517}),
    .b({net_150,net_452}),
    .c({net_151,open_n97}),
    .d({net_228,net_1141}),
    .mi({io_mcu_d[1],io_mcu_d[0]}),
    .f({net_238,net_235}),
    .q({net_229,net_228})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hC0C0"),
    .INIT_LUTG0("16'hC8C8"),
    .INIT_LUTF1("16'hA0A0"),
    .INIT_LUTG1("16'hA0A0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_177
  (
    .a({net_316,net_249}),
    .b({open_n98,i_mcu_rws}),
    .c({i_mcu_rws,i_mcu_dcs}),
    .e({open_n99,net_316}),
    .f({net_236,net_234})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hAF23"),
    .INIT_LUTG0("16'h0A02"),
    .INIT_LUTF1("16'h0501"),
    .INIT_LUTG1("16'h5511"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_178
  (
    .clk(gclk_9),
    .ce(net_304),
    .a({net_232,net_230}),
    .b({net_302,net_178}),
    .c({net_231,net_233}),
    .d({net_163,net_231}),
    .e({net_178,net_144}),
    .mi({io_mcu_d[1],io_mcu_d[0]}),
    .f({net_237,net_232}),
    .q({net_231,net_230})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_179
  (
    .clk(gclk_5),
    .sr(net_90),
    .mi({open_n100,net_170}),
    .q({open_n101,net_233})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hE000"),
    .INIT_LUT1("16'hCCC8"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_180
  (
    .clk(gclk_5),
    .sr(net_90),
    .a({net_1141,net_239}),
    .b({net_1349,net_155}),
    .c({net_1283,net_163}),
    .d({net_324,net_176}),
    .mi({open_n102,net_157}),
    .f({net_241,net_240}),
    .q({open_n103,net_239})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h4F04"),
    .INIT_LUTG0("16'hFF0F"),
    .INIT_LUTF1("16'h00F5"),
    .INIT_LUTG1("16'hF5F5"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_181
  (
    .clk(gclk_9),
    .ce(net_304),
    .a({net_243,net_242}),
    .b({open_n104,net_87}),
    .c({net_88,net_303}),
    .d({net_242,net_174}),
    .e({net_87,net_307}),
    .mi({io_mcu_d[5],io_mcu_d[6]}),
    .f({net_245,net_246}),
    .q({net_243,net_242})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h030A"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_182
  (
    .a({net_85,net_85}),
    .b({net_252,net_252}),
    .c({net_181,net_181}),
    .d({net_180,net_180}),
    .mi({open_n105,net_896}),
    .fx({open_n106,net_244})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h5F3F"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_183
  (
    .a({net_723,net_723}),
    .b({net_716,net_716}),
    .c({net_1044,net_189}),
    .d({net_189,net_1044}),
    .mi({open_n107,net_186}),
    .fx({open_n108,net_250})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h8AAA"),
    .INIT_LUTG0("16'hBAAA"),
    .INIT_LUTF1("16'hFAAA"),
    .INIT_LUTG1("16'h8AAA"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_184
  (
    .clk(gclk_9),
    .ce(net_184),
    .a({net_248,net_247}),
    .b({net_180,net_181}),
    .c({net_647,net_308}),
    .d({net_308,net_647}),
    .e({net_181,net_180}),
    .q({net_248,net_247})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'hA000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h4444"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_185
  (
    .clk(gclk_9),
    .ce(net_251),
    .a({net_180,net_308}),
    .b({net_181,open_n109}),
    .c({open_n110,net_181}),
    .d({open_n111,net_180}),
    .e({net_308,net_895}),
    .mi({open_n112,io_mcu_d[0]}),
    .f({net_249,net_251}),
    .q({open_n113,net_253})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h5F3F"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_186
  (
    .a({net_721,net_721}),
    .b({net_715,net_715}),
    .c({net_189,net_189}),
    .d({net_1044,net_1044}),
    .mi({open_n114,net_258}),
    .fx({open_n115,net_252})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0100"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_187
  (
    .a({net_321,net_321}),
    .b({net_260,net_260}),
    .c({net_338,net_338}),
    .d({net_1114,net_1114}),
    .mi({open_n116,net_244}),
    .fx({open_n117,net_254})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hCC55"),
    .INIT_LUTG0("16'hF0F0"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h50F0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_188
  (
    .clk(gclk_9),
    .a({net_1341,net_257}),
    .b({open_n118,net_530}),
    .c({net_814,net_256}),
    .d({net_256,i_mcu_dcs}),
    .e({net_466,i_mcu_rws}),
    .f({net_257,open_n119}),
    .q({open_n120,net_256})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h00A0"),
    .INIT_LUTG0("16'h00A0"),
    .INIT_LUTF1("16'hAA00"),
    .INIT_LUTG1("16'hAA00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_189
  (
    .clk(gclk_8),
    .ce(net_261),
    .sr(net_182),
    .a({net_648,net_564}),
    .c({open_n121,net_847}),
    .d({net_255,net_247}),
    .mi({open_n122,io_i2c_sda}),
    .f({net_260,net_261}),
    .q({open_n123,net_255})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0A0C"),
    .INIT_LUT1("16'h0503"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_190
  (
    .a({net_61,net_733}),
    .b({net_51,net_743}),
    .c({net_189,net_189}),
    .d({net_1044,net_1044}),
    .f({net_259,net_258})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'hCCCC"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hFF00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_191
  (
    .b({open_n124,net_998}),
    .d({i_mcu_rws,open_n125}),
    .e({net_547,i_mcu_rws}),
    .f({net_265,net_264})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h888A"),
    .INIT_LUTG0("16'h88FA"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h57DF"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_192
  (
    .clk(gclk_9),
    .a({net_959,net_263}),
    .b({net_1301,net_793}),
    .c({net_196,net_264}),
    .d({net_263,i_mcu_dcs}),
    .e({net_197,io_mcu_d[5]}),
    .f({net_266,open_n126}),
    .q({open_n127,net_263})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hCC0F"),
    .INIT_LUT1("16'hFF00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_193
  (
    .clk(gclk_9),
    .a({net_559,net_262}),
    .b({net_643,net_643}),
    .c({i_mcu_dcs,net_559}),
    .d({net_262,i_mcu_dcs}),
    .mi({open_n128,i_mcu_rws}),
    .q({open_n129,net_262})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h888A"),
    .INIT_LUTG0("16'h8F8A"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hDD55"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_194
  (
    .clk(gclk_9),
    .a({net_199,net_267}),
    .b({net_592,net_793}),
    .c({open_n130,i_mcu_dcs}),
    .d({net_267,net_264}),
    .e({net_1523,io_mcu_d[1]}),
    .f({net_269,open_n131}),
    .q({open_n132,net_267})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hBBAA"),
    .INIT_LUTG0("16'hBBB0"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hEAC0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_195
  (
    .clk(gclk_9),
    .a({net_943,net_268}),
    .b({net_277,net_793}),
    .c({net_1155,io_mcu_d[6]}),
    .d({net_268,i_mcu_dcs}),
    .e({net_950,net_100}),
    .f({net_270,open_n133}),
    .q({open_n134,net_268})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h0700"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_196
  (
    .a({net_968,net_968}),
    .b({net_205,net_205}),
    .c({net_345,net_345}),
    .d({net_204,net_204}),
    .mi({open_n135,net_498}),
    .fx({open_n136,net_276})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h7F0F"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0B00"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_197
  (
    .a({net_488,net_585}),
    .b({net_862,net_101}),
    .c({net_273,net_961}),
    .d({net_272,net_209}),
    .e({net_270,net_203}),
    .f({net_274,net_272})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h888A"),
    .INIT_LUTG0("16'h8F8A"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hEAC0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_198
  (
    .clk(gclk_9),
    .a({net_964,net_271}),
    .b({net_104,net_793}),
    .c({net_961,i_mcu_dcs}),
    .d({net_271,net_265}),
    .e({net_592,io_mcu_d[4]}),
    .f({net_273,open_n137}),
    .q({open_n138,net_271})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0A00"),
    .INIT_LUT1("16'hFF0B"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_199
  (
    .clk(gclk_9),
    .a({io_mcu_d[3],io_mcu_d[3]}),
    .b({net_265,net_793}),
    .c({i_mcu_dcs,i_mcu_dcs}),
    .d({net_793,net_265}),
    .mi({open_n139,net_275}),
    .q({open_n140,net_275})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hBBAA"),
    .INIT_LUT1("16'hFC54"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_200
  (
    .clk(gclk_9),
    .a({net_793,net_277}),
    .b({io_mcu_d[5],net_793}),
    .c({i_mcu_dcs,io_mcu_d[5]}),
    .d({net_277,i_mcu_dcs}),
    .mi({open_n141,net_343}),
    .q({open_n142,net_277})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hBBAA"),
    .INIT_LUTG0("16'hBBB0"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hDD55"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_201
  (
    .clk(gclk_9),
    .a({net_213,net_278}),
    .b({net_1521,net_793}),
    .c({open_n143,io_mcu_d[2]}),
    .d({net_278,i_mcu_dcs}),
    .e({net_962,net_343}),
    .f({net_281,open_n144}),
    .q({open_n145,net_278})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h888A"),
    .INIT_LUTG0("16'h8F8A"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hEAC0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_202
  (
    .clk(gclk_9),
    .a({net_951,net_279}),
    .b({net_215,net_793}),
    .c({net_564,i_mcu_dcs}),
    .d({net_279,net_265}),
    .e({net_863,io_mcu_d[0]}),
    .f({net_282,open_n146}),
    .q({open_n147,net_279})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0A00"),
    .INIT_LUT1("16'hCECF"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_203
  (
    .clk(gclk_9),
    .a({io_mcu_d[6],io_mcu_d[6]}),
    .b({net_793,net_793}),
    .c({i_mcu_dcs,i_mcu_dcs}),
    .d({net_344,net_344}),
    .mi({open_n148,net_280}),
    .q({open_n149,net_280})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hF000"),
    .INIT_LUT1("16'h0F0F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_204
  (
    .c({i_mcu_rws,i_mcu_rws}),
    .d({open_n150,net_1113}),
    .f({net_288,net_286})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h888A"),
    .INIT_LUTG0("16'h88FA"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hECA0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_205
  (
    .clk(gclk_9),
    .a({net_862,net_284}),
    .b({net_952,net_793}),
    .c({net_289,net_286}),
    .d({net_284,i_mcu_dcs}),
    .e({net_668,io_mcu_d[0]}),
    .f({net_287,open_n151}),
    .q({open_n152,net_284})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h888A"),
    .INIT_LUTG0("16'h8F8A"),
    .INIT_LUTF1("16'h888A"),
    .INIT_LUTG1("16'h8F8A"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_206
  (
    .clk(gclk_9),
    .a({net_283,net_285}),
    .b({net_793,net_793}),
    .c({i_mcu_dcs,i_mcu_dcs}),
    .d({net_286,net_286}),
    .e({io_mcu_d[4],io_mcu_d[7]}),
    .q({net_283,net_285})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0808"),
    .INIT_LUT1("16'hFF0B"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_207
  (
    .clk(gclk_9),
    .a({io_mcu_d[3],io_mcu_d[3]}),
    .b({net_286,net_286}),
    .c({i_mcu_dcs,i_mcu_dcs}),
    .d({net_793,net_793}),
    .mi({open_n153,net_289}),
    .q({open_n154,net_289})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hCE0A"),
    .INIT_LUT1("16'hCE0A"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_212
  (
    .clk(gclk_9),
    .a({net_290,net_291}),
    .b({net_109,net_125}),
    .c({net_234,net_234}),
    .d({net_512,net_512}),
    .q({net_290,net_291})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_213
  (
    .clk(gclk_0),
    .sr(net_451),
    .mi({net_395,net_392}),
    .q({net_292,net_293})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_214
  (
    .clk(gclk_0),
    .sr(net_451),
    .mi({net_413,net_382}),
    .q({net_297,net_294})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_215
  (
    .clk(gclk_0),
    .sr(net_451),
    .mi({net_391,net_390}),
    .q({net_295,net_296})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_216
  (
    .clk(gclk_0),
    .sr(net_451),
    .mi({net_410,net_426}),
    .q({net_298,net_299})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hAF23"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hAA00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_217
  (
    .clk(gclk_9),
    .ce(net_304),
    .a({net_1283,net_301}),
    .b({open_n155,net_163}),
    .c({open_n156,net_162}),
    .d({net_452,net_302}),
    .e({net_517,net_237}),
    .mi({io_mcu_d[2],io_mcu_d[3]}),
    .f({net_304,net_305}),
    .q({net_302,net_301})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'hD0DD"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h50DC"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_218
  (
    .clk(gclk_9),
    .ce(net_304),
    .a({net_300,net_303}),
    .b({net_88,net_174}),
    .c({net_166,net_166}),
    .d({net_243,net_300}),
    .e({net_245,net_245}),
    .mi({io_mcu_d[4],io_mcu_d[7]}),
    .f({net_307,net_306}),
    .q({net_300,net_303})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h2222"),
    .INIT_LUTG0("16'h2222"),
    .INIT_LUTF1("16'h0003"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_219
  (
    .a({open_n157,net_644}),
    .b({net_530,net_643}),
    .c({net_314,open_n158}),
    .d({net_645,open_n159}),
    .e({net_531,open_n160}),
    .f({net_309,net_308})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hCC00"),
    .INIT_LUT1("16'h4545"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_220
  (
    .clk(gclk_9),
    .ce(net_313),
    .a({net_1341,open_n161}),
    .b({net_1141,net_1141}),
    .c({net_916,open_n162}),
    .d({open_n163,net_446}),
    .mi({open_n164,io_mcu_d[0]}),
    .f({net_310,net_313}),
    .q({open_n165,net_311})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h0100"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_221
  (
    .a({net_181,net_181}),
    .b({net_644,net_644}),
    .c({net_643,net_643}),
    .d({net_180,net_180}),
    .mi({open_n166,net_316}),
    .fx({open_n167,net_312})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h1100"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0004"),
    .INIT_LUTG1("16'h0004"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_222
  (
    .clk(gclk_9),
    .ce(net_184),
    .a({net_530,net_314}),
    .b({net_531,net_531}),
    .c({net_645,open_n168}),
    .d({net_314,net_645}),
    .e({open_n169,net_530}),
    .mi({open_n170,io_mcu_d[7]}),
    .f({net_316,net_315}),
    .q({open_n171,net_314})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0500"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h00CC"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_223
  (
    .clk(gclk_9),
    .ce(net_320),
    .a({open_n172,net_181}),
    .b({net_180,open_n173}),
    .c({open_n174,net_180}),
    .d({net_181,net_308}),
    .e({net_308,net_895}),
    .mi({open_n175,io_mcu_d[0]}),
    .f({net_319,net_320}),
    .q({open_n176,net_322})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hBB00"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0B00"),
    .INIT_LUTG1("16'h0B00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_224
  (
    .clk(gclk_9),
    .ce(net_454),
    .a({net_317,net_318}),
    .b({net_1283,net_1283}),
    .c({net_331,open_n177}),
    .d({net_312,net_312}),
    .e({open_n178,net_328}),
    .mi({io_mcu_d[7],io_mcu_d[3]}),
    .f({net_321,net_323}),
    .q({net_317,net_318})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hCC0F"),
    .INIT_LUT1("16'hFF00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_225
  (
    .clk(gclk_9),
    .a({net_807,net_324}),
    .b({net_645,net_645}),
    .c({i_mcu_dcs,net_807}),
    .d({net_324,i_mcu_dcs}),
    .mi({open_n179,i_mcu_rws}),
    .q({open_n180,net_324})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h1133"),
    .INIT_LUTG0("16'h1100"),
    .INIT_LUTF1("16'h0033"),
    .INIT_LUTG1("16'h1111"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_226
  (
    .clk(gclk_9),
    .ce(net_535),
    .a({net_326,net_325}),
    .b({net_1283,net_1283}),
    .d({net_190,net_1141}),
    .e({net_1141,net_262}),
    .mi({io_mcu_d[6],io_mcu_d[3]}),
    .f({net_327,net_328}),
    .q({net_326,net_325})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h5F3F"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_227
  (
    .a({net_717,net_717}),
    .b({net_711,net_711}),
    .c({net_189,net_189}),
    .d({net_1044,net_1044}),
    .mi({open_n181,net_183}),
    .fx({open_n182,net_329})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0503"),
    .INIT_LUTG0("16'h0503"),
    .INIT_LUTF1("16'h4400"),
    .INIT_LUTG1("16'hCC88"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_228
  (
    .clk(gclk_9),
    .ce(net_535),
    .a({net_1141,net_330}),
    .b({net_439,net_188}),
    .c({open_n183,net_1283}),
    .d({net_188,net_1141}),
    .e({net_1150,open_n184}),
    .mi({open_n185,io_mcu_d[7]}),
    .f({net_332,net_331}),
    .q({open_n186,net_330})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h00A0"),
    .INIT_LUT1("16'hF000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_229
  (
    .clk(gclk_8),
    .ce(net_337),
    .sr(net_182),
    .a({open_n187,net_1056}),
    .c({net_1113,net_668}),
    .d({net_333,net_247}),
    .mi({open_n188,io_i2c_sda}),
    .f({net_338,net_337}),
    .q({open_n189,net_333})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h8888"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'hC0C0"),
    .INIT_LUTG1("16'hEEEE"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_230
  (
    .clk(gclk_8),
    .ce(net_340),
    .sr(net_182),
    .a({net_1276,net_1276}),
    .b({net_1067,net_668}),
    .c({net_1468,open_n190}),
    .e({net_951,net_247}),
    .mi({open_n191,io_i2c_sda}),
    .f({net_334,net_340}),
    .q({open_n192,net_336})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hB000"),
    .INIT_LUT1("16'h00AA"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_231
  (
    .a({net_1038,net_310}),
    .b({open_n193,net_188}),
    .c({open_n194,net_554}),
    .d({net_266,net_254}),
    .f({net_335,net_339})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hFFFF"),
    .INIT_LUT1("16'hDF0F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("INV"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_232
  (
    .clk(gclk_8),
    .ce(net_248),
    .a({net_1532,net_341}),
    .b({net_487,net_1532}),
    .c({net_574,net_487}),
    .d({net_341,net_574}),
    .mi({open_n195,net_680}),
    .q({open_n196,net_341})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'hF0F0"),
    .INIT_LUTF1("16'hA0A0"),
    .INIT_LUTG1("16'hA0A0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_233
  (
    .a({net_906,open_n197}),
    .c({i_mcu_rws,i_mcu_rws}),
    .e({open_n198,net_999}),
    .f({net_344,net_343})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h2FAF"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("INV"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_234
  (
    .clk(gclk_8),
    .ce(net_248),
    .a({net_489,net_342}),
    .b({net_346,net_346}),
    .c({net_481,net_481}),
    .d({net_342,net_489}),
    .mi({open_n199,net_582}),
    .q({open_n200,net_342})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'hA000"),
    .INIT_LUTF1("16'h0022"),
    .INIT_LUTG1("16'h2222"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_235
  (
    .a({net_350,net_1289}),
    .b({net_826,open_n201}),
    .c({open_n202,net_962}),
    .d({net_849,net_202}),
    .e({net_962,net_960}),
    .f({net_346,net_345})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h01FF"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_236
  (
    .a({net_843,net_843}),
    .b({net_668,net_952}),
    .c({net_862,net_862}),
    .d({net_952,net_668}),
    .mi({open_n203,net_477}),
    .fx({open_n204,net_348})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0007"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h8000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_237
  (
    .a({net_347,net_352}),
    .b({net_485,net_207}),
    .c({net_361,net_355}),
    .d({net_509,net_335}),
    .e({net_276,net_281}),
    .f({net_349,net_347})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h1000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_238
  (
    .a({net_968,net_475}),
    .b({net_475,net_968}),
    .c({net_572,net_572}),
    .d({net_570,net_570}),
    .mi({open_n205,net_860}),
    .fx({open_n206,net_350})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hA000"),
    .INIT_LUT1("16'h8888"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_239
  (
    .a({net_951,net_843}),
    .b({net_952,open_n207}),
    .c({open_n208,net_275}),
    .d({open_n209,net_951}),
    .f({net_352,net_355})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h888A"),
    .INIT_LUTG0("16'h8F8A"),
    .INIT_LUTF1("16'hA000"),
    .INIT_LUTG1("16'hA000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_240
  (
    .clk(gclk_9),
    .a({net_843,net_351}),
    .b({open_n210,net_793}),
    .c({net_1032,i_mcu_dcs}),
    .d({net_351,net_344}),
    .e({open_n211,io_mcu_d[4]}),
    .f({net_353,open_n212}),
    .q({open_n213,net_351})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h001F"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_241
  (
    .a({net_950,net_950}),
    .b({net_862,net_862}),
    .c({net_951,net_951}),
    .d({net_588,net_588}),
    .mi({open_n214,net_840}),
    .fx({open_n215,net_354})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hBBAA"),
    .INIT_LUTG0("16'hBBB0"),
    .INIT_LUTF1("16'h8800"),
    .INIT_LUTG1("16'h8800"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_242
  (
    .clk(gclk_9),
    .a({net_951,net_356}),
    .b({net_950,net_793}),
    .c({open_n216,io_mcu_d[2]}),
    .d({net_356,i_mcu_dcs}),
    .e({open_n217,net_265}),
    .f({net_357,open_n218}),
    .q({open_n219,net_356})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hBBAA"),
    .INIT_LUTG0("16'hBBB0"),
    .INIT_LUTF1("16'hF000"),
    .INIT_LUTG1("16'hF000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_243
  (
    .clk(gclk_9),
    .a({open_n220,net_358}),
    .b({open_n221,net_793}),
    .c({net_475,io_mcu_d[7]}),
    .d({net_358,i_mcu_dcs}),
    .e({open_n222,net_343}),
    .f({net_359,open_n223}),
    .q({open_n224,net_358})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0A00"),
    .INIT_LUT1("16'hCECF"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_244
  (
    .clk(gclk_9),
    .a({io_mcu_d[6],io_mcu_d[6]}),
    .b({net_793,net_793}),
    .c({i_mcu_dcs,i_mcu_dcs}),
    .d({net_286,net_286}),
    .mi({open_n225,net_360}),
    .q({open_n226,net_360})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0001"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_245
  (
    .a({net_359,net_359}),
    .b({net_579,net_579}),
    .c({net_590,net_590}),
    .d({net_595,net_595}),
    .mi({open_n227,net_282}),
    .fx({open_n228,net_361})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0A00"),
    .INIT_LUT1("16'hAEAF"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_246
  (
    .clk(gclk_9),
    .a({net_793,io_mcu_d[5]}),
    .b({io_mcu_d[5],net_793}),
    .c({i_mcu_dcs,i_mcu_dcs}),
    .d({net_344,net_344}),
    .mi({open_n229,net_364}),
    .q({open_n230,net_364})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h888A"),
    .INIT_LUTG0("16'h8F8A"),
    .INIT_LUTF1("16'h8A8A"),
    .INIT_LUTG1("16'h8F88"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_247
  (
    .clk(gclk_9),
    .a({net_363,net_362}),
    .b({net_793,net_793}),
    .c({i_mcu_dcs,i_mcu_dcs}),
    .d({io_mcu_d[3],net_344}),
    .e({net_344,io_mcu_d[2]}),
    .q({net_363,net_362})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h000A"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB_CARRY"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_248
  (
    .clk(gclk_0),
    .sr(net_451),
    .a({net_635,open_n231}),
    .b({net_377,open_n232}),
    .mi({net_378,net_379}),
    .q({net_368,net_366}),
    .fco(block_248_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_249
  (
    .clk(gclk_9),
    .ce(net_634),
    .a({net_365,net_367}),
    .b({net_366,net_374}),
    .mi({io_mcu_d[2],io_mcu_d[1]}),
    .fci(block_248_carry),
    .q({net_365,net_367}),
    .fco(block_249_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_250
  (
    .clk(gclk_9),
    .ce(net_634),
    .a({net_370,net_372}),
    .b({net_380,net_373}),
    .mi({io_mcu_d[4],io_mcu_d[3]}),
    .fci(block_249_carry),
    .q({net_370,net_372}),
    .fco(block_250_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_251
  (
    .clk(gclk_9),
    .ce(net_634),
    .a({net_369,net_371}),
    .b({net_294,net_368}),
    .mi({io_mcu_d[6],io_mcu_d[5]}),
    .fci(block_250_carry),
    .q({net_369,net_371}),
    .fco(block_251_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_252
  (
    .clk(gclk_9),
    .ce(net_634),
    .a({net_1130,net_376}),
    .b({net_293,net_400}),
    .mi({open_n233,io_mcu_d[7]}),
    .fci(block_251_carry),
    .q({open_n234,net_376}),
    .fco(block_252_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_255
  (
    .clk(gclk_9),
    .ce(net_640),
    .a({net_639,net_375}),
    .b({net_389,net_296}),
    .mi({open_n235,io_mcu_d[1]}),
    .fci(block_252_carry),
    .q({open_n236,net_375}),
    .fco(block_255_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_256
  (
    .clk(gclk_9),
    .ce(net_640),
    .a({net_396,net_638}),
    .b({net_399,net_387}),
    .mi({open_n237,io_mcu_d[4]}),
    .fci(block_255_carry),
    .q({open_n238,net_396}),
    .fco(block_256_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_259
  (
    .clk(gclk_9),
    .ce(net_640),
    .a({net_386,net_388}),
    .b({net_292,net_295}),
    .mi({io_mcu_d[6],io_mcu_d[5]}),
    .fci(block_256_carry),
    .q({net_386,net_388}),
    .fco(block_259_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_260
  (
    .clk(gclk_9),
    .ce(net_640),
    .a({net_311,net_405}),
    .b({net_411,net_401}),
    .mi({open_n239,io_mcu_d[7]}),
    .fci(block_259_carry),
    .q({open_n240,net_405}),
    .fco(block_260_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_263
  (
    .clk(gclk_9),
    .ce(net_313),
    .a({net_402,net_404}),
    .b({net_521,net_297}),
    .mi({io_mcu_d[2],io_mcu_d[1]}),
    .fci(block_260_carry),
    .q({net_402,net_404}),
    .fco(block_263_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_264
  (
    .clk(gclk_9),
    .ce(net_313),
    .a({net_418,net_421}),
    .b({net_407,net_403}),
    .mi({io_mcu_d[4],io_mcu_d[3]}),
    .fci(block_263_carry),
    .q({net_418,net_421}),
    .fco(block_264_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_267
  (
    .clk(gclk_9),
    .ce(net_313),
    .a({net_417,net_420}),
    .b({net_298,net_520}),
    .mi({io_mcu_d[6],io_mcu_d[5]}),
    .fci(block_264_carry),
    .q({net_417,net_420}),
    .fco(block_267_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_268
  (
    .clk(gclk_9),
    .ce(net_313),
    .a({net_456,net_435}),
    .b({net_427,net_416}),
    .mi({open_n241,io_mcu_d[7]}),
    .fci(block_267_carry),
    .q({open_n242,net_435}),
    .fco(block_268_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_270
  (
    .clk(gclk_9),
    .ce(net_455),
    .a({net_433,net_434}),
    .b({net_518,net_299}),
    .mi({io_mcu_d[2],io_mcu_d[1]}),
    .fci(block_268_carry),
    .q({net_433,net_434}),
    .fco(block_270_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_272
  (
    .clk(gclk_9),
    .ce(net_455),
    .a({net_441,net_443}),
    .b({net_422,net_419}),
    .mi({io_mcu_d[4],io_mcu_d[3]}),
    .fci(block_270_carry),
    .q({net_441,net_443}),
    .fco(block_272_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_274
  (
    .clk(gclk_9),
    .ce(net_455),
    .a({net_440,net_442}),
    .b({net_522,net_438}),
    .mi({io_mcu_d[6],io_mcu_d[5]}),
    .fci(block_272_carry),
    .q({net_440,net_442}),
    .fco(block_274_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_276
  (
    .clk(gclk_9),
    .ce(net_455),
    .a({1'b0,net_450}),
    .b({open_n243,net_432}),
    .mi({open_n244,io_mcu_d[7]}),
    .fci(block_274_carry),
    .f({net_451,open_n245}),
    .q({open_n246,net_450})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h000A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_253
  (
    .clk(gclk_0),
    .sr(net_451),
    .a({net_374,1'b0}),
    .b({net_366,net_377}),
    .c({1'b0,1'b0}),
    .d({1'b0,open_n247}),
    .e({1'b0,open_n248}),
    .mi({net_381,net_385}),
    .f({net_381,open_n249}),
    .fx({net_379,net_385}),
    .q({net_374,net_377}),
    .fco(sig_253_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_254
  (
    .clk(gclk_0),
    .sr(net_451),
    .a({net_368,net_373}),
    .b({net_294,net_380}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_383,net_384}),
    .fci(sig_253_carry),
    .f({net_378,net_384}),
    .fx({net_382,net_383}),
    .q({net_380,net_373}),
    .fco(sig_254_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_257
  (
    .clk(gclk_0),
    .sr(net_451),
    .a({net_296,net_400}),
    .b({net_389,net_293}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_394,net_398}),
    .fci(sig_254_carry),
    .f({net_390,net_394}),
    .fx({net_398,net_392}),
    .q({net_400,net_389}),
    .fco(sig_257_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_258
  (
    .clk(gclk_0),
    .sr(net_451),
    .a({net_295,net_387}),
    .b({net_292,net_399}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_393,net_397}),
    .fci(sig_257_carry),
    .f({net_391,net_397}),
    .fx({net_395,net_393}),
    .q({net_399,net_387}),
    .fco(sig_258_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_261
  (
    .clk(gclk_0),
    .sr(net_451),
    .a({net_297,net_401}),
    .b({net_521,net_411}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_414,net_409}),
    .fci(sig_258_carry),
    .f({net_413,net_409}),
    .fx({net_408,net_414}),
    .q({net_411,net_401}),
    .fco(sig_261_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_262
  (
    .clk(gclk_0),
    .sr(net_451),
    .a({net_520,net_403}),
    .b({net_298,net_407}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_412,net_415}),
    .fci(sig_261_carry),
    .f({net_406,net_415}),
    .fx({net_410,net_412}),
    .q({net_407,net_403}),
    .fco(sig_262_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_265
  (
    .clk(gclk_0),
    .sr(net_451),
    .a({net_299,net_416}),
    .b({net_518,net_427}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_429,net_424}),
    .fci(sig_262_carry),
    .f({net_426,net_424}),
    .fx({net_423,net_429}),
    .q({net_427,net_416}),
    .fco(sig_265_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_266
  (
    .clk(gclk_0),
    .sr(net_451),
    .a({net_438,net_419}),
    .b({net_522,net_422}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_428,net_431}),
    .fci(sig_265_carry),
    .f({net_430,net_431}),
    .fx({net_425,net_428}),
    .q({net_422,net_419}),
    .fco(sig_266_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_269
  (
    .clk(gclk_0),
    .sr(net_451),
    .a({open_n250,net_432}),
    .c({1'b0,1'b0}),
    .d({open_n251,1'b0}),
    .mi({net_430,net_437}),
    .fci(sig_266_carry),
    .f({open_n252,net_437}),
    .q({net_438,net_432})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h8080"),
    .INIT_LUTF1("16'h1000"),
    .INIT_LUTG1("16'h1000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_271
  (
    .a({net_181,net_308}),
    .b({net_180,net_647}),
    .c({net_308,net_181}),
    .d({net_315,open_n253}),
    .e({open_n254,net_180}),
    .f({net_439,net_436})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h00BF"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'hF33F"),
    .INIT_LUTG1("16'h033F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_273
  (
    .clk(gclk_9),
    .ce(net_535),
    .a({open_n255,net_444}),
    .b({net_309,net_644}),
    .c({net_181,net_643}),
    .d({net_180,net_220}),
    .e({net_647,net_532}),
    .mi({open_n256,io_mcu_d[5]}),
    .f({net_444,net_447}),
    .q({open_n257,net_448})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0100"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h4000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_275
  (
    .clk(gclk_9),
    .ce(net_449),
    .a({net_181,net_181}),
    .b({net_224,net_644}),
    .c({net_180,net_643}),
    .d({net_644,net_180}),
    .e({net_643,net_224}),
    .mi({open_n258,io_mcu_d[0]}),
    .f({net_446,net_449}),
    .q({open_n259,net_445})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h00CC"),
    .INIT_LUTG0("16'h00CC"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h8888"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_277
  (
    .clk(gclk_9),
    .ce(net_454),
    .a({net_452,open_n260}),
    .b({net_532,i_mcu_rws}),
    .d({open_n261,i_mcu_dcs}),
    .e({net_1283,open_n262}),
    .mi({io_mcu_d[2],io_mcu_d[1]}),
    .f({net_454,net_452}),
    .q({net_457,net_458})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hAA00"),
    .INIT_LUT1("16'hAA00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_278
  (
    .clk(gclk_9),
    .ce(net_455),
    .a({net_525,net_1283}),
    .d({net_1283,net_446}),
    .mi({open_n263,io_mcu_d[0]}),
    .f({net_453,net_455}),
    .q({open_n264,net_456})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0BBB"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_279
  (
    .a({net_250,net_250}),
    .b({net_523,net_523}),
    .c({net_1113,net_1113}),
    .d({net_336,net_336}),
    .mi({open_n265,net_653}),
    .fx({open_n266,net_467})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hF0CC"),
    .INIT_LUTG0("16'hAAAA"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h0777"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_280
  (
    .clk(gclk_9),
    .ce(net_454),
    .a({net_547,net_460}),
    .b({net_471,net_256}),
    .c({net_312,net_448}),
    .d({net_462,net_1141}),
    .e({net_1238,net_1283}),
    .mi({open_n267,io_mcu_d[5]}),
    .f({net_466,net_462}),
    .q({open_n268,net_460})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0503"),
    .INIT_LUT1("16'h4404"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_281
  (
    .clk(gclk_9),
    .ce(net_535),
    .a({net_464,net_461}),
    .b({net_312,net_908}),
    .c({net_1283,net_1283}),
    .d({net_457,net_1141}),
    .mi({open_n269,io_mcu_d[2]}),
    .f({net_465,net_464}),
    .q({open_n270,net_461})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0080"),
    .INIT_LUTF1("16'hA0F0"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_282
  (
    .clk(gclk_9),
    .ce(net_454),
    .a({net_459,net_931}),
    .b({open_n271,net_467}),
    .c({net_312,net_659}),
    .d({net_1283,net_463}),
    .e({net_327,net_1505}),
    .mi({io_mcu_d[6],open_n272}),
    .f({net_463,net_468}),
    .q({net_459,open_n273})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h5000"),
    .INIT_LUT1("16'h050F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_283
  (
    .clk(gclk_8),
    .ce(net_473),
    .sr(net_182),
    .a({net_906,net_247}),
    .c({net_332,net_1032}),
    .d({net_469,net_1067}),
    .mi({open_n274,io_i2c_sda}),
    .f({net_472,net_473}),
    .q({open_n275,net_469})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA0A0"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h8888"),
    .INIT_LUTG1("16'h8888"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_284
  (
    .clk(gclk_8),
    .ce(net_474),
    .sr(net_182),
    .a({net_1056,net_1056}),
    .b({net_1289,open_n276}),
    .c({open_n277,net_951}),
    .e({open_n278,net_247}),
    .mi({open_n279,io_i2c_sda}),
    .f({net_470,net_474}),
    .q({open_n280,net_471})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0088"),
    .INIT_LUT1("16'hC0C0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_285
  (
    .clk(gclk_8),
    .ce(net_479),
    .sr(net_182),
    .a({open_n281,net_1056}),
    .b({net_1468,net_1468}),
    .c({net_950,open_n282}),
    .d({open_n283,net_247}),
    .mi({open_n284,io_i2c_sda}),
    .f({net_475,net_479}),
    .q({open_n285,net_482})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h4040"),
    .INIT_LUTG0("16'h4040"),
    .INIT_LUTF1("16'hF0C0"),
    .INIT_LUTG1("16'hF0F0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_286
  (
    .clk(gclk_8),
    .ce(net_476),
    .sr(net_182),
    .a({open_n286,net_247}),
    .b({net_1276,net_847}),
    .c({net_1032,net_1032}),
    .d({net_843,open_n287}),
    .e({net_863,open_n288}),
    .mi({open_n289,io_i2c_sda}),
    .f({net_477,net_476}),
    .q({open_n290,net_478})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h00A0"),
    .INIT_LUTG0("16'h00A0"),
    .INIT_LUTF1("16'h7777"),
    .INIT_LUTG1("16'h0077"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_287
  (
    .clk(gclk_8),
    .ce(net_483),
    .sr(net_182),
    .a({net_564,net_847}),
    .b({net_847,open_n291}),
    .c({open_n292,net_951}),
    .d({net_1523,net_247}),
    .e({net_862,open_n293}),
    .mi({open_n294,io_i2c_sda}),
    .f({net_480,net_483}),
    .q({open_n295,net_484})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h035F"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_288
  (
    .a({net_1060,net_1060}),
    .b({net_863,net_863}),
    .c({net_952,net_952}),
    .d({net_584,net_584}),
    .mi({open_n296,net_247}),
    .fx({open_n297,net_481})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h0001"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_289
  (
    .a({net_269,net_269}),
    .b({net_493,net_493}),
    .c({net_1245,net_1245}),
    .d({net_353,net_353}),
    .mi({open_n298,net_494}),
    .fx({open_n299,net_485})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h4040"),
    .INIT_LUTF1("16'h8888"),
    .INIT_LUTG1("16'h8888"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_290
  (
    .a({net_570,net_487}),
    .b({net_580,net_497}),
    .c({open_n300,net_575}),
    .e({open_n301,net_672}),
    .f({net_487,net_489})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hBBAA"),
    .INIT_LUTG0("16'hBBB0"),
    .INIT_LUTF1("16'h3333"),
    .INIT_LUTG1("16'h0033"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_291
  (
    .clk(gclk_9),
    .a({open_n302,net_486}),
    .b({net_967,net_793}),
    .c({open_n303,io_mcu_d[0]}),
    .d({net_486,i_mcu_dcs}),
    .e({net_961,net_816}),
    .f({net_488,open_n304}),
    .q({open_n305,net_486})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h0007"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_292
  (
    .a({net_1060,net_1060}),
    .b({net_1067,net_1067}),
    .c({net_969,net_969}),
    .d({net_588,net_588}),
    .mi({open_n306,net_838}),
    .fx({open_n307,net_490})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0D00"),
    .INIT_LUT1("16'h0500"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_293
  (
    .a({net_674,net_668}),
    .b({open_n308,net_211}),
    .c({net_334,net_357}),
    .d({net_958,net_502}),
    .f({net_497,net_498})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h001F"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h1000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_294
  (
    .a({net_688,net_962}),
    .b({net_1068,net_863}),
    .c({net_354,net_668}),
    .d({net_492,net_968}),
    .e({net_348,net_826}),
    .f({net_495,net_492})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h888A"),
    .INIT_LUTG0("16'h8F8A"),
    .INIT_LUTF1("16'h050F"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_295
  (
    .clk(gclk_9),
    .a({net_969,net_491}),
    .b({open_n309,net_793}),
    .c({net_593,i_mcu_dcs}),
    .d({net_491,net_344}),
    .e({net_287,io_mcu_d[7]}),
    .f({net_494,open_n310}),
    .q({open_n311,net_491})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h8800"),
    .INIT_LUT1("16'h2222"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_296
  (
    .a({net_668,net_283}),
    .b({net_1067,net_950}),
    .d({open_n312,net_668}),
    .f({net_496,net_493})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0777"),
    .INIT_LUT1("16'hA0A0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_297
  (
    .a({net_1468,net_1523}),
    .b({open_n313,net_950}),
    .c({net_585,net_843}),
    .d({open_n314,net_1468}),
    .f({net_499,net_500})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hBBAA"),
    .INIT_LUTG0("16'hBBB0"),
    .INIT_LUTF1("16'h7F7F"),
    .INIT_LUTG1("16'h007F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_298
  (
    .clk(gclk_9),
    .a({net_285,net_501}),
    .b({net_843,net_793}),
    .c({net_1333,io_mcu_d[1]}),
    .d({net_501,i_mcu_dcs}),
    .e({net_499,net_100}),
    .f({net_503,open_n315}),
    .q({open_n316,net_501})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h7F0F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_299
  (
    .a({net_863,net_863}),
    .b({net_508,net_508}),
    .c({net_1521,net_1521}),
    .d({net_594,net_594}),
    .mi({open_n317,net_247}),
    .fx({open_n318,net_502})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0A00"),
    .INIT_LUT1("16'hCECF"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_300
  (
    .clk(gclk_9),
    .a({io_mcu_d[3],io_mcu_d[3]}),
    .b({net_793,net_793}),
    .c({i_mcu_dcs,i_mcu_dcs}),
    .d({net_343,net_343}),
    .mi({open_n319,net_508}),
    .q({open_n320,net_508})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hBBAA"),
    .INIT_LUTG0("16'hBBB0"),
    .INIT_LUTF1("16'h8080"),
    .INIT_LUTG1("16'hAA80"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_301
  (
    .clk(gclk_9),
    .a({net_1032,net_505}),
    .b({net_950,net_793}),
    .c({net_363,io_mcu_d[1]}),
    .d({net_505,i_mcu_dcs}),
    .e({net_863,net_344}),
    .f({net_507,open_n321}),
    .q({open_n322,net_505})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hBBAA"),
    .INIT_LUTG0("16'hBBB0"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h0111"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_302
  (
    .clk(gclk_9),
    .a({net_685,net_506}),
    .b({net_507,net_793}),
    .c({net_684,io_mcu_d[0]}),
    .d({net_506,i_mcu_dcs}),
    .e({net_503,net_100}),
    .f({net_509,open_n323}),
    .q({open_n324,net_506})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hBBAA"),
    .INIT_LUT1("16'hFC54"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_303
  (
    .clk(gclk_9),
    .a({net_793,net_504}),
    .b({i_mcu_dcs,net_793}),
    .c({io_mcu_d[7],io_mcu_d[7]}),
    .d({net_504,i_mcu_dcs}),
    .mi({open_n325,net_100}),
    .q({open_n326,net_504})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hF000"),
    .INIT_LUT1("16'h0808"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_304
  (
    .clk(gclk_9),
    .ce(net_513),
    .a({net_249,open_n327}),
    .b({net_236,open_n328}),
    .c({i_mcu_dcs,net_222}),
    .d({open_n329,net_249}),
    .mi({open_n330,io_mcu_d[0]}),
    .f({net_512,net_513}),
    .q({open_n331,net_511})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0100"),
    .INIT_LUTF1("16'h00F0"),
    .INIT_LUTG1("16'hFFF0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_305
  (
    .clk(gclk_9),
    .ce(net_515),
    .a({open_n332,i_mcu_dcs}),
    .b({open_n333,net_180}),
    .c({gclk_2,net_181}),
    .d({net_510,net_1111}),
    .e({net_1337,net_236}),
    .mi({open_n334,io_mcu_d[0]}),
    .f({net_514,net_515}),
    .q({open_n335,net_510})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hC0C0"),
    .INIT_LUTG0("16'hC0C0"),
    .INIT_LUTF1("16'hF000"),
    .INIT_LUTG1("16'hF000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_306
  (
    .clk(gclk_9),
    .ce(net_519),
    .b({open_n336,net_222}),
    .c({net_319,net_319}),
    .d({net_533,open_n337}),
    .mi({open_n338,io_mcu_d[0]}),
    .f({net_517,net_519}),
    .q({open_n339,net_516})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_307
  (
    .clk(gclk_0),
    .sr(net_451),
    .mi({net_406,net_423}),
    .q({net_520,net_518})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_308
  (
    .clk(gclk_0),
    .sr(net_451),
    .mi({net_408,net_425}),
    .q({net_521,net_522})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h8000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_309
  (
    .a({net_315,net_315}),
    .b({net_180,net_180}),
    .c({net_181,net_181}),
    .d({net_644,net_644}),
    .mi({open_n340,net_643}),
    .fx({open_n341,net_525})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h8000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h0100"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_310
  (
    .clk(gclk_9),
    .ce(net_526),
    .a({net_180,net_224}),
    .b({net_644,net_180}),
    .c({net_643,net_181}),
    .d({net_533,net_644}),
    .e({net_181,net_643}),
    .mi({open_n342,io_mcu_d[0]}),
    .f({net_524,net_526}),
    .q({open_n343,net_527})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h00F0"),
    .INIT_LUTF1("16'h2222"),
    .INIT_LUTG1("16'h2222"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_311
  (
    .a({net_523,open_n344}),
    .b({net_528,open_n345}),
    .c({open_n346,net_896}),
    .d({open_n347,net_181}),
    .e({open_n348,net_180}),
    .f({net_529,net_523})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h5F3F"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_312
  (
    .a({net_720,net_720}),
    .b({net_708,net_708}),
    .c({net_189,net_189}),
    .d({net_1044,net_1044}),
    .mi({open_n349,net_666}),
    .fx({open_n350,net_528})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0002"),
    .INIT_LUT1("16'h0400"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_313
  (
    .clk(gclk_9),
    .ce(net_184),
    .a({net_531,net_530}),
    .b({net_645,net_645}),
    .c({net_314,net_314}),
    .d({net_530,net_531}),
    .mi({io_mcu_d[6],io_mcu_d[5]}),
    .f({net_533,net_536}),
    .q({net_531,net_530})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0400"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hF000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_314
  (
    .clk(gclk_9),
    .ce(net_535),
    .a({open_n351,net_180}),
    .b({open_n352,net_533}),
    .c({net_1141,net_181}),
    .d({net_532,net_644}),
    .e({net_452,net_643}),
    .mi({io_mcu_d[0],io_mcu_d[4]}),
    .f({net_535,net_532}),
    .q({net_538,net_534})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0777"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_315
  (
    .a({net_905,net_905}),
    .b({net_642,net_642}),
    .c({net_648,net_648}),
    .d({net_482,net_482}),
    .mi({open_n353,net_637}),
    .fx({open_n354,net_537})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0088"),
    .INIT_LUTG0("16'h0088"),
    .INIT_LUTF1("16'h0FFF"),
    .INIT_LUTG1("16'h0555"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_316
  (
    .clk(gclk_8),
    .ce(net_541),
    .sr(net_182),
    .a({net_874,net_1468}),
    .b({open_n355,net_1067}),
    .c({net_648,open_n356}),
    .d({net_539,net_247}),
    .e({net_905,open_n357}),
    .mi({open_n358,io_i2c_sda}),
    .f({net_540,net_541}),
    .q({open_n359,net_539})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hF0CC"),
    .INIT_LUTG0("16'hAAAA"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h0777"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_317
  (
    .clk(gclk_9),
    .ce(net_454),
    .a({net_1341,net_543}),
    .b({net_324,net_324}),
    .c({net_312,net_534}),
    .d({net_545,net_1141}),
    .e({net_1049,net_1283}),
    .mi({open_n360,io_mcu_d[4]}),
    .f({net_548,net_545}),
    .q({open_n361,net_543})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h5050"),
    .INIT_LUTG0("16'h5050"),
    .INIT_LUTF1("16'hCC00"),
    .INIT_LUTG1("16'hCC00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_318
  (
    .clk(gclk_8),
    .ce(net_550),
    .sr(net_182),
    .a({open_n362,net_247}),
    .b({net_1113,open_n363}),
    .c({open_n364,net_957}),
    .d({net_544,open_n365}),
    .mi({open_n366,io_i2c_sda}),
    .f({net_546,net_550}),
    .q({open_n367,net_544})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h2020"),
    .INIT_LUT1("16'h020A"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_319
  (
    .clk(gclk_8),
    .ce(net_549),
    .sr(net_182),
    .a({net_540,net_1161}),
    .b({net_1113,net_247}),
    .c({net_633,net_1303}),
    .d({net_542,open_n368}),
    .mi({open_n369,io_i2c_sda}),
    .f({net_551,net_549}),
    .q({open_n370,net_542})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h4000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_320
  (
    .a({net_181,net_181}),
    .b({net_180,net_180}),
    .c({net_647,net_647}),
    .d({net_644,net_644}),
    .mi({open_n371,net_643}),
    .fx({open_n372,net_547})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h2020"),
    .INIT_LUT1("16'h0BBB"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_321
  (
    .clk(gclk_8),
    .ce(net_556),
    .sr(net_182),
    .a({net_651,net_847}),
    .b({net_523,net_247}),
    .c({net_1113,net_668}),
    .d({net_552,open_n373}),
    .mi({open_n374,io_i2c_sda}),
    .f({net_557,net_556}),
    .q({open_n375,net_552})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0C00"),
    .INIT_LUTG0("16'h0C00"),
    .INIT_LUTF1("16'hC0C0"),
    .INIT_LUTG1("16'h00C0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_322
  (
    .clk(gclk_8),
    .ce(net_555),
    .sr(net_182),
    .b({net_1108,net_1648}),
    .c({net_472,net_247}),
    .d({net_553,net_1528}),
    .e({net_547,open_n376}),
    .mi({open_n377,io_i2c_sda}),
    .f({net_554,net_555}),
    .q({open_n378,net_553})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0777"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h8A8A"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_323
  (
    .a({net_558,net_547}),
    .b({net_310,net_484}),
    .c({net_262,net_1053}),
    .d({open_n379,net_906}),
    .e({net_795,net_1515}),
    .f({net_559,net_558})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h00A0"),
    .INIT_LUT1("16'h153F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_324
  (
    .clk(gclk_8),
    .ce(net_566),
    .sr(net_182),
    .a({net_547,net_951}),
    .b({net_478,open_n380}),
    .c({net_906,net_1276}),
    .d({net_560,net_247}),
    .mi({open_n381,io_i2c_sda}),
    .f({net_565,net_566}),
    .q({open_n382,net_560})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0444"),
    .INIT_LUTG0("16'h0404"),
    .INIT_LUTF1("16'hEEC0"),
    .INIT_LUTG1("16'hEEC0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_325
  (
    .a({net_847,net_562}),
    .b({net_1276,net_561}),
    .c({net_1521,net_1161}),
    .d({net_1468,net_470}),
    .e({open_n383,net_1528}),
    .f({net_562,net_563})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0777"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h0888"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_326
  (
    .a({net_561,net_1333}),
    .b({net_571,net_1276}),
    .c({net_1525,net_1056}),
    .d({net_1047,net_1468}),
    .e({net_348,net_957}),
    .f({net_567,net_561})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hE000"),
    .INIT_LUT1("16'hAA00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_327
  (
    .a({net_943,net_961}),
    .b({open_n384,net_943}),
    .c({open_n385,net_847}),
    .d({net_1289,net_1289}),
    .f({net_564,net_568})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0FFF"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h00CC"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_328
  (
    .b({net_567,open_n386}),
    .c({open_n387,net_1528}),
    .d({net_829,net_1648}),
    .e({net_836,net_352}),
    .f({net_570,net_571})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h1000"),
    .INIT_LUT1("16'h1000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_329
  (
    .a({net_968,net_1068}),
    .b({net_475,net_1161}),
    .c({net_490,net_681}),
    .d({net_846,net_480}),
    .f({net_569,net_572})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h5554"),
    .INIT_LUTF1("16'h0005"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_330
  (
    .a({net_1047,net_687}),
    .b({open_n388,net_961}),
    .c({net_670,net_1302}),
    .d({net_1303,net_573}),
    .e({net_1528,net_848}),
    .f({net_573,net_574})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h8000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_331
  (
    .a({net_489,net_489}),
    .b({net_860,net_860}),
    .c({net_495,net_495}),
    .d({net_563,net_563}),
    .mi({open_n389,net_686}),
    .fx({open_n390,net_578})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0777"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h8000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_332
  (
    .a({net_495,net_564}),
    .b({net_497,net_950}),
    .c({net_682,net_1155}),
    .d({net_575,net_853}),
    .e({net_850,net_499}),
    .f({net_580,net_575})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0700"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h333B"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_333
  (
    .a({net_576,net_966}),
    .b({net_342,net_1329}),
    .c({net_487,net_851}),
    .d({net_1065,net_682}),
    .e({net_349,net_852}),
    .f({net_582,net_576})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0088"),
    .INIT_LUT1("16'h2F00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_334
  (
    .clk(gclk_8),
    .ce(net_581),
    .sr(net_182),
    .a({net_1525,net_1525}),
    .b({net_586,net_1303}),
    .c({net_274,open_n391}),
    .d({net_1289,net_247}),
    .mi({open_n392,io_i2c_sda}),
    .f({net_579,net_581}),
    .q({open_n393,net_577})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hC0C0"),
    .INIT_LUT1("16'hAA00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_335
  (
    .a({net_584,open_n394}),
    .b({open_n395,net_961}),
    .c({open_n396,net_1289}),
    .d({net_962,open_n397}),
    .f({net_588,net_584})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hBBAA"),
    .INIT_LUTG0("16'hBBB0"),
    .INIT_LUTF1("16'h030F"),
    .INIT_LUTG1("16'h0105"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_336
  (
    .clk(gclk_9),
    .a({net_862,net_583}),
    .b({net_962,net_793}),
    .c({net_587,io_mcu_d[0]}),
    .d({net_583,i_mcu_dcs}),
    .e({net_362,net_344}),
    .f({net_586,open_n398}),
    .q({open_n399,net_583})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hAC00"),
    .INIT_LUT1("16'h2222"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_337
  (
    .a({net_1078,net_364}),
    .b({net_1301,net_280}),
    .c({open_n400,net_1301}),
    .d({open_n401,net_1078}),
    .f({net_585,net_587})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h888A"),
    .INIT_LUTG0("16'h8F8A"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hAA00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_338
  (
    .clk(gclk_9),
    .a({net_585,net_589}),
    .b({open_n402,net_793}),
    .c({open_n403,i_mcu_dcs}),
    .d({net_589,net_343}),
    .e({net_1333,io_mcu_d[0]}),
    .f({net_590,open_n404}),
    .q({open_n405,net_589})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'hCCCC"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hCC00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_339
  (
    .b({net_668,net_1078}),
    .d({net_592,open_n406}),
    .e({net_360,net_1301}),
    .f({net_593,net_592})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h888A"),
    .INIT_LUTG0("16'h8F8A"),
    .INIT_LUTF1("16'h153F"),
    .INIT_LUTG1("16'h153F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_340
  (
    .clk(gclk_9),
    .a({net_952,net_591}),
    .b({net_843,net_793}),
    .c({net_596,i_mcu_dcs}),
    .d({net_591,net_343}),
    .e({open_n407,io_mcu_d[1]}),
    .f({net_594,open_n408}),
    .q({open_n409,net_591})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'hF888"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_341
  (
    .a({net_1523,net_1523}),
    .b({net_504,net_504}),
    .c({net_1521,net_1521}),
    .d({net_597,net_597}),
    .mi({open_n410,net_862}),
    .fx({open_n411,net_595})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h888A"),
    .INIT_LUTG0("16'h8F8A"),
    .INIT_LUTF1("16'hBBAA"),
    .INIT_LUTG1("16'hBBB0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_342
  (
    .clk(gclk_9),
    .a({net_597,net_596}),
    .b({net_793,net_793}),
    .c({io_mcu_d[4],i_mcu_dcs}),
    .d({i_mcu_dcs,net_343}),
    .e({net_343,io_mcu_d[6]}),
    .q({net_597,net_596})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0B0B"),
    .INIT_LUTG0("16'h0B00"),
    .INIT_LUTF1("16'hC4F5"),
    .INIT_LUTG1("16'hC4F5"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_347
  (
    .clk(gclk_9),
    .ce(net_612),
    .a({net_599,net_598}),
    .b({net_745,net_752}),
    .c({net_775,net_601}),
    .d({net_610,net_599}),
    .e({open_n412,net_775}),
    .mi({io_mcu_d[5],io_mcu_d[4]}),
    .f({net_604,net_606}),
    .q({net_599,net_598})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hAF23"),
    .INIT_LUTG0("16'h0A02"),
    .INIT_LUTF1("16'h0501"),
    .INIT_LUTG1("16'h5511"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_348
  (
    .clk(gclk_9),
    .ce(net_612),
    .a({net_603,net_600}),
    .b({net_602,net_747}),
    .c({net_598,net_615}),
    .d({net_747,net_602}),
    .e({net_752,net_773}),
    .mi({io_mcu_d[3],io_mcu_d[2]}),
    .f({net_601,net_603}),
    .q({net_602,net_600})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_349
  (
    .clk(gclk_5),
    .sr(net_880),
    .mi({open_n413,net_763}),
    .q({open_n414,net_605})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h5D04"),
    .INIT_LUTG0("16'hFF55"),
    .INIT_LUTF1("16'h5050"),
    .INIT_LUTG1("16'h5050"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_350
  (
    .clk(gclk_9),
    .ce(net_612),
    .a({net_610,net_608}),
    .b({open_n415,net_604}),
    .c({net_745,net_606}),
    .d({open_n416,net_767}),
    .e({open_n417,net_613}),
    .mi({io_mcu_d[6],io_mcu_d[7]}),
    .f({net_613,net_611}),
    .q({net_610,net_608})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h8888"),
    .INIT_LUTF1("16'h50F5"),
    .INIT_LUTG1("16'hF5F5"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_351
  (
    .clk(gclk_9),
    .ce(net_612),
    .a({net_607,net_524}),
    .b({open_n418,net_1141}),
    .c({net_748,open_n419}),
    .d({net_609,open_n420}),
    .e({net_749,net_452}),
    .mi({io_mcu_d[1],io_mcu_d[0]}),
    .f({net_615,net_612}),
    .q({net_607,net_609})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h5F3F"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_352
  (
    .a({net_705,net_705}),
    .b({net_697,net_697}),
    .c({net_1044,net_904}),
    .d({net_904,net_1044}),
    .mi({open_n421,net_189}),
    .fx({open_n422,net_614})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h000A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD_CARRY"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("F"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_353
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_617,1'b0}),
    .q({net_617,open_n423}),
    .fco(block_353_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_354
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_616,net_618}),
    .b({1'b0,1'b0}),
    .fci(block_353_carry),
    .q({net_616,net_618}),
    .fco(block_354_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_355
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({open_n424,net_620}),
    .b({open_n425,1'b0}),
    .fci(block_354_carry),
    .q({open_n426,net_620})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h7777"),
    .INIT_LUTG0("16'h2222"),
    .INIT_LUTF1("16'h3333"),
    .INIT_LUTG1("16'h0F0F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_356
  (
    .a({open_n427,net_516}),
    .b({net_85,net_873}),
    .c({net_1212,open_n428}),
    .e({net_516,net_147}),
    .f({net_623,net_624})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hAF23"),
    .INIT_LUTG0("16'h0A02"),
    .INIT_LUTF1("16'h1101"),
    .INIT_LUTG1("16'h5505"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_357
  (
    .clk(gclk_9),
    .ce(net_779),
    .a({net_622,net_619}),
    .b({net_777,net_744}),
    .c({net_621,net_611}),
    .d({net_744,net_621}),
    .e({net_761,net_605}),
    .mi({io_mcu_d[1],io_mcu_d[0]}),
    .f({net_625,net_622}),
    .q({net_621,net_619})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h0C0A"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_358
  (
    .a({net_147,net_147}),
    .b({net_873,net_873}),
    .c({net_180,net_180}),
    .d({net_181,net_181}),
    .mi({open_n429,net_896}),
    .fx({open_n430,net_626})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h1000"),
    .INIT_LUT1("16'h0F55"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_359
  (
    .a({net_146,net_180}),
    .b({open_n431,net_181}),
    .c({net_874,net_146}),
    .d({net_516,net_896}),
    .f({net_630,net_633})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h2020"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h5555"),
    .INIT_LUTG1("16'h00FF"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_360
  (
    .a({net_161,net_896}),
    .b({open_n432,net_181}),
    .c({open_n433,net_161}),
    .d({net_1083,open_n434}),
    .e({net_516,net_180}),
    .f({net_631,net_628})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hFEFA"),
    .INIT_LUT1("16'h11DD"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_361
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_709,net_627}),
    .b({net_1044,net_616}),
    .c({open_n435,net_620}),
    .d({net_719,net_618}),
    .f({net_629,open_n436}),
    .q({open_n437,net_627})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h1000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h0101"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_362
  (
    .clk(gclk_9),
    .ce(net_634),
    .a({net_524,net_1264}),
    .b({net_517,net_1508}),
    .c({net_525,net_1263}),
    .d({open_n438,net_446}),
    .e({net_447,net_1507}),
    .mi({open_n439,io_mcu_d[0]}),
    .f({net_632,net_634}),
    .q({open_n440,net_635})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h1000"),
    .INIT_LUT1("16'h05F5"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_363
  (
    .a({net_86,net_180}),
    .b({open_n441,net_181}),
    .c({net_516,net_86}),
    .d({net_642,net_896}),
    .f({net_636,net_637})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0001"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h0004"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_364
  (
    .clk(gclk_9),
    .ce(net_640),
    .a({net_1507,io_mcu_d[7]}),
    .b({net_446,io_mcu_d[6]}),
    .c({net_1264,io_mcu_d[5]}),
    .d({net_1508,io_mcu_d[4]}),
    .e({net_1263,io_mcu_d[3]}),
    .mi({io_mcu_d[2],io_mcu_d[3]}),
    .f({net_640,net_641}),
    .q({net_639,net_638})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hAFCF"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_365
  (
    .a({net_722,net_722}),
    .b({net_712,net_712}),
    .c({net_189,net_189}),
    .d({net_1044,net_1044}),
    .mi({open_n442,net_664}),
    .fx({open_n443,net_642})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h4000"),
    .INIT_LUT1("16'h0008"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_366
  (
    .a({net_315,net_181}),
    .b({net_1111,net_180}),
    .c({net_181,net_647}),
    .d({net_180,net_1111}),
    .f({net_652,net_648})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'hF5FF"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h0404"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_367
  (
    .clk(gclk_9),
    .ce(net_184),
    .a({net_645,net_643}),
    .b({net_531,open_n444}),
    .c({net_314,net_181}),
    .d({open_n445,net_647}),
    .e({net_530,net_1010}),
    .mi({io_mcu_d[4],io_mcu_d[3]}),
    .f({net_647,net_649}),
    .q({net_645,net_643})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h1008"),
    .INIT_LUTF1("16'h0040"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_368
  (
    .clk(gclk_9),
    .ce(net_184),
    .a({net_646,net_644}),
    .b({net_911,net_180}),
    .c({net_1341,net_643}),
    .d({net_436,net_181}),
    .e({net_652,net_309}),
    .mi({open_n446,io_mcu_d[2]}),
    .f({net_650,net_646}),
    .q({open_n447,net_644})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h5F3F"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_369
  (
    .a({net_724,net_724}),
    .b({net_713,net_713}),
    .c({net_189,net_189}),
    .d({net_1044,net_1044}),
    .mi({open_n448,net_657}),
    .fx({open_n449,net_651})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'hC00A"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_370
  (
    .a({net_179,net_179}),
    .b({net_1555,net_1555}),
    .c({net_180,net_180}),
    .d({net_181,net_181}),
    .mi({open_n450,net_896}),
    .fx({open_n451,net_653})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0404"),
    .INIT_LUTG0("16'h5454"),
    .INIT_LUTF1("16'h2233"),
    .INIT_LUTG1("16'h0011"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_371
  (
    .a({net_1044,net_189}),
    .b({net_189,net_742}),
    .c({open_n452,net_1044}),
    .d({net_741,open_n453}),
    .e({net_732,net_731}),
    .f({net_658,net_657})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hFF4F"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0311"),
    .INIT_LUTG1("16'h0311"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_372
  (
    .clk(gclk_4),
    .ce(net_1291),
    .sr(net_445),
    .a({net_262,net_655}),
    .b({net_1283,net_1283}),
    .c({net_927,net_439}),
    .d({net_1141,net_656}),
    .e({open_n454,net_323}),
    .mi({open_n455,net_1288}),
    .f({net_656,net_661}),
    .q({open_n456,net_655})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h2020"),
    .INIT_LUT1("16'h0777"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_373
  (
    .clk(gclk_8),
    .ce(net_660),
    .sr(net_182),
    .a({net_905,net_670}),
    .b({net_987,net_247}),
    .c({net_648,net_943}),
    .d({net_654,open_n457}),
    .mi({open_n458,io_i2c_sda}),
    .f({net_659,net_660}),
    .q({open_n459,net_654})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0A0C"),
    .INIT_LUT1("16'h0053"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_374
  (
    .a({net_728,net_729}),
    .b({net_738,net_737}),
    .c({net_1044,net_189}),
    .d({net_189,net_1044}),
    .f({net_664,net_666})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hCC55"),
    .INIT_LUTG0("16'hF0F0"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h44CC"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_375
  (
    .clk(gclk_9),
    .a({net_1341,net_663}),
    .b({net_810,net_181}),
    .c({open_n460,net_662}),
    .d({net_662,i_mcu_dcs}),
    .e({net_803,i_mcu_rws}),
    .f({net_663,open_n461}),
    .q({open_n462,net_662})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0FFF"),
    .INIT_LUT1("16'h0111"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_376
  (
    .a({net_662,net_662}),
    .b({net_1141,net_1141}),
    .c({net_669,net_669}),
    .d({net_1113,net_1113}),
    .mi({open_n463,net_916}),
    .fx({open_n464,net_665})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hA0A0"),
    .INIT_LUT1("16'hF000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_377
  (
    .clk(gclk_8),
    .ce(net_667),
    .sr(net_182),
    .a({open_n465,net_920}),
    .c({net_1161,net_1161}),
    .d({net_1289,open_n466}),
    .mi({open_n467,io_i2c_sda}),
    .f({net_668,net_667}),
    .q({open_n468,net_669})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h3030"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hCCCC"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_378
  (
    .clk(gclk_8),
    .ce(net_673),
    .sr(net_182),
    .b({net_1289,net_247}),
    .c({open_n469,net_951}),
    .e({net_929,net_929}),
    .mi({open_n470,io_i2c_sda}),
    .f({net_670,net_673}),
    .q({open_n471,net_671})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0070"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_379
  (
    .a({net_1333,net_1333}),
    .b({net_1067,net_1067}),
    .c({net_841,net_841}),
    .d({net_829,net_829}),
    .mi({open_n472,net_949}),
    .fx({open_n473,net_672})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h00C0"),
    .INIT_LUT1("16'hF8A8"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_380
  (
    .clk(gclk_8),
    .ce(net_675),
    .sr(net_182),
    .a({net_1521,open_n474}),
    .b({net_1299,net_929}),
    .c({net_843,net_1521}),
    .d({net_951,net_247}),
    .mi({open_n475,io_i2c_sda}),
    .f({net_674,net_675}),
    .q({open_n476,net_676})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hBBBB"),
    .INIT_LUT1("16'h000B"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_381
  (
    .a({net_1532,net_1532}),
    .b({net_1057,net_1057}),
    .c({net_670,net_1047}),
    .d({net_1047,net_670}),
    .mi({open_n477,net_961}),
    .fx({open_n478,net_677})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h8000"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h5000"),
    .INIT_LUTG1("16'h5500"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_382
  (
    .a({net_965,net_679}),
    .b({open_n479,net_563}),
    .c({net_1532,net_677}),
    .d({net_854,net_955}),
    .e({net_857,net_334}),
    .f({net_679,net_680})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0777"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h22AA"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_383
  (
    .a({net_678,net_584}),
    .b({net_951,net_863}),
    .c({open_n480,net_1032}),
    .d({net_962,net_952}),
    .e({net_500,net_965}),
    .f({net_682,net_678})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h007F"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_384
  (
    .a({net_851,net_470}),
    .b({net_470,net_963}),
    .c({net_963,net_1302}),
    .d({net_1302,net_851}),
    .mi({open_n481,net_969}),
    .fx({open_n482,net_681})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hFFFE"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_385
  (
    .a({net_496,net_496}),
    .b({net_1068,net_1032}),
    .c({net_1032,net_1068}),
    .d({net_970,net_970}),
    .mi({open_n483,net_1532}),
    .fx({open_n484,net_687})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0505"),
    .INIT_LUTG0("16'h4444"),
    .INIT_LUTF1("16'hF000"),
    .INIT_LUTG1("16'hF000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_386
  (
    .a({open_n485,net_684}),
    .b({open_n486,net_1532}),
    .c({net_1468,net_964}),
    .d({net_592,open_n487}),
    .e({open_n488,net_1300}),
    .f({net_684,net_686})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h888A"),
    .INIT_LUTG0("16'h8F8A"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hF888"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_387
  (
    .clk(gclk_9),
    .a({net_964,net_683}),
    .b({net_689,net_793}),
    .c({net_1648,i_mcu_dcs}),
    .d({net_683,net_265}),
    .e({net_966,io_mcu_d[7]}),
    .f({net_685,open_n489}),
    .q({open_n490,net_683})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hB000"),
    .INIT_LUT1("16'hCCCC"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_388
  (
    .a({net_1532,net_1300}),
    .b({net_1060,net_1532}),
    .c({net_1301,net_1301}),
    .d({net_1300,net_1060}),
    .mi({open_n491,net_1299}),
    .fx({open_n492,net_688})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0A00"),
    .INIT_LUT1("16'hFF0B"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_389
  (
    .clk(gclk_9),
    .a({io_mcu_d[5],io_mcu_d[5]}),
    .b({net_265,net_793}),
    .c({i_mcu_dcs,i_mcu_dcs}),
    .d({net_793,net_265}),
    .mi({open_n493,net_689}),
    .q({open_n494,net_689})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_411
  (
    .clk(gclk_5),
    .sr(net_880),
    .mi({net_755,net_764}),
    .q({net_745,net_744})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hCCAA"),
    .INIT_LUT1("16'h0F0F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_412
  (
    .clk(gclk_4),
    .a({net_759,net_746}),
    .b({net_994,net_759}),
    .c({net_511,net_511}),
    .d({net_746,net_994}),
    .mi({open_n495,net_445}),
    .q({open_n496,net_746})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h000A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_413
  (
    .clk(gclk_5),
    .sr(net_880),
    .a({net_748,1'b0}),
    .b({net_773,net_749}),
    .c({1'b0,1'b0}),
    .d({1'b0,open_n497}),
    .e({1'b0,open_n498}),
    .mi({net_753,net_758}),
    .f({net_753,open_n499}),
    .fx({net_751,net_758}),
    .q({net_748,net_749}),
    .fco(sig_413_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_414
  (
    .clk(gclk_5),
    .sr(net_880),
    .a({net_775,net_747}),
    .b({net_745,net_752}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_754,net_757}),
    .fci(sig_413_carry),
    .f({net_756,net_757}),
    .fx({net_755,net_754}),
    .q({net_752,net_747}),
    .fco(sig_414_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_416
  (
    .clk(gclk_5),
    .sr(net_880),
    .a({net_744,net_767}),
    .b({net_761,net_605}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_768,net_771}),
    .fci(sig_414_carry),
    .f({net_764,net_768}),
    .fx({net_771,net_763}),
    .q({net_767,net_761}),
    .fco(sig_416_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_417
  (
    .clk(gclk_5),
    .sr(net_880),
    .a({net_878,net_760}),
    .b({net_877,net_762}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_765,net_770}),
    .fci(sig_416_carry),
    .f({net_769,net_770}),
    .fx({net_766,net_765}),
    .q({net_762,net_760}),
    .fco(sig_417_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_419
  (
    .clk(gclk_5),
    .sr(net_880),
    .a({open_n500,net_772}),
    .c({1'b0,1'b0}),
    .d({open_n501,1'b0}),
    .mi({net_751,net_774}),
    .fci(sig_417_carry),
    .f({open_n502,net_774}),
    .q({net_773,net_772})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h5F3F"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_415
  (
    .a({net_702,net_702}),
    .b({net_690,net_690}),
    .c({net_1044,net_904}),
    .d({net_904,net_1044}),
    .mi({open_n503,net_189}),
    .fx({open_n504,net_750})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h33AA"),
    .INIT_LUT1("16'h3333"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_418
  (
    .clk(gclk_4),
    .a({net_636,net_759}),
    .b({net_511,net_636}),
    .c({net_994,net_511}),
    .d({net_759,net_994}),
    .mi({open_n505,net_445}),
    .q({open_n506,net_759})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'hEFFF"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_420
  (
    .a({net_181,net_181}),
    .b({net_180,net_180}),
    .c({net_896,net_896}),
    .d({net_160,net_160}),
    .mi({open_n507,net_786}),
    .fx({open_n508,net_780})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'hE0E0"),
    .INIT_LUTF1("16'h0101"),
    .INIT_LUTG1("16'h0101"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_421
  (
    .clk(gclk_5),
    .sr(net_880),
    .a({net_439,net_775}),
    .b({net_312,net_752}),
    .c({net_1349,net_761}),
    .e({open_n509,net_745}),
    .mi({open_n510,net_756}),
    .f({net_778,net_782}),
    .q({open_n511,net_775})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hAF23"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hF000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_422
  (
    .clk(gclk_9),
    .ce(net_779),
    .a({open_n512,net_776}),
    .b({open_n513,net_761}),
    .c({net_1283,net_760}),
    .d({net_524,net_777}),
    .e({net_452,net_625}),
    .mi({io_mcu_d[2],io_mcu_d[3]}),
    .f({net_779,net_784}),
    .q({net_777,net_776})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h1B1B"),
    .INIT_LUT1("16'h4747"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_423
  (
    .a({net_787,net_516}),
    .b({net_516,net_95}),
    .c({net_160,net_1209}),
    .f({net_781,net_783})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h7F7F"),
    .INIT_LUT1("16'h1555"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_424
  (
    .a({net_436,net_319}),
    .b({net_309,net_309}),
    .c({net_627,net_627}),
    .d({net_319,net_436}),
    .mi({open_n514,net_1062}),
    .fx({open_n515,net_786})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hF4FF"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'hE000"),
    .INIT_LUTG1("16'hF000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("INV"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_425
  (
    .clk(gclk_5),
    .ce(net_90),
    .a({net_1005,net_162}),
    .b({net_1002,net_301}),
    .c({net_1009,net_305}),
    .d({net_1001,net_306}),
    .e({net_1003,net_246}),
    .f({net_785,open_n516}),
    .q({open_n517,net_788})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hAFCF"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_426
  (
    .a({net_725,net_725}),
    .b({net_714,net_714}),
    .c({net_189,net_189}),
    .d({net_1044,net_1044}),
    .mi({open_n518,net_658}),
    .fx({open_n519,net_787})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hBB0B"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h020A"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_427
  (
    .a({net_789,net_985}),
    .b({net_652,net_904}),
    .c({net_918,net_523}),
    .d({net_1348,net_91}),
    .e({net_804,net_546}),
    .f({net_790,net_789})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h1000"),
    .INIT_LUTF1("16'h8888"),
    .INIT_LUTG1("16'h8888"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_428
  (
    .a({net_905,net_792}),
    .b({net_1083,net_529}),
    .c({open_n520,net_797}),
    .d({open_n521,net_661}),
    .e({open_n522,net_913}),
    .f({net_792,net_795})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hFF00"),
    .INIT_LUTG0("16'h5F00"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hFF00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_429
  (
    .clk(gclk_4),
    .a({open_n523,net_647}),
    .c({open_n524,i_mcu_rws}),
    .d({net_536,i_mcu_dcs}),
    .e({net_319,net_319}),
    .mi({i_adc1A_d[3],open_n525}),
    .f({net_794,net_793}),
    .q({net_799,open_n526})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0808"),
    .INIT_LUT1("16'h020A"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_430
  (
    .clk(gclk_8),
    .ce(net_798),
    .sr(net_182),
    .a({net_1345,net_1047}),
    .b({net_1113,net_1161}),
    .c({net_628,net_247}),
    .d({net_791,open_n527}),
    .mi({open_n528,io_i2c_sda}),
    .f({net_797,net_798}),
    .q({open_n529,net_791})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h4000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_431
  (
    .a({net_180,net_180}),
    .b({net_647,net_647}),
    .c({net_181,net_181}),
    .d({net_644,net_644}),
    .mi({open_n530,net_643}),
    .fx({open_n531,net_796})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h4040"),
    .INIT_LUT1("16'h0777"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_432
  (
    .clk(gclk_8),
    .ce(net_805),
    .sr(net_182),
    .a({net_905,net_247}),
    .b({net_787,net_1276}),
    .c({net_648,net_1468}),
    .d({net_800,open_n532}),
    .mi({open_n533,io_i2c_sda}),
    .f({net_804,net_805}),
    .q({open_n534,net_800})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0777"),
    .INIT_LUTF1("16'h8000"),
    .INIT_LUTG1("16'h8000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_433
  (
    .clk(gclk_4),
    .a({net_665,net_1251}),
    .b({net_947,i_adc2A_d[1]}),
    .c({net_537,net_796}),
    .d({net_802,net_932}),
    .e({open_n535,net_1518}),
    .mi({open_n536,i_adc2A_d[1]}),
    .f({net_803,net_802}),
    .q({open_n537,net_806})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hB000"),
    .INIT_LUT1("16'h8000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_434
  (
    .a({net_565,net_181}),
    .b({net_915,net_1041}),
    .c({net_1121,net_548}),
    .d({net_1491,net_801}),
    .f({net_801,net_807})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hAACC"),
    .INIT_LUTG0("16'hF0F0"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h153F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_435
  (
    .clk(gclk_9),
    .ce(net_535),
    .a({net_809,net_808}),
    .b({net_439,net_662}),
    .c({net_1160,net_458}),
    .d({net_312,net_1141}),
    .e({net_993,net_1283}),
    .mi({open_n538,io_mcu_d[1]}),
    .f({net_810,net_809}),
    .q({open_n539,net_808})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0777"),
    .INIT_LUT1("16'h8888"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_436
  (
    .clk(gclk_4),
    .a({i_mcu_rws,net_796}),
    .b({net_796,net_828}),
    .c({open_n540,i_adc1A_d[7]}),
    .d({open_n541,net_1244}),
    .mi({open_n542,i_adc1A_d[7]}),
    .f({net_816,net_820}),
    .q({open_n543,net_819})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0777"),
    .INIT_LUTF1("16'h0400"),
    .INIT_LUTG1("16'h0400"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_437
  (
    .clk(gclk_4),
    .a({net_1030,net_794}),
    .b({net_813,i_adc1B_d[5]}),
    .c({net_626,net_796}),
    .d({net_811,net_941}),
    .e({open_n544,net_936}),
    .mi({open_n545,i_adc1B_d[5]}),
    .f({net_814,net_811}),
    .q({open_n546,net_818})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0777"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h4444"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_438
  (
    .clk(gclk_8),
    .ce(net_817),
    .sr(net_182),
    .a({net_247,net_904}),
    .b({net_943,net_1556}),
    .c({open_n547,net_648}),
    .d({open_n548,net_812}),
    .e({net_1047,net_557}),
    .mi({io_i2c_sda,open_n549}),
    .f({net_817,net_813}),
    .q({net_812,open_n550})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0777"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_439
  (
    .a({net_547,net_547}),
    .b({net_671,net_671}),
    .c({net_1527,net_1527}),
    .d({net_906,net_906}),
    .mi({open_n551,net_465}),
    .fx({open_n552,net_815})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h4040"),
    .INIT_LUT1("16'h8888"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_440
  (
    .clk(gclk_8),
    .ce(net_825),
    .sr(net_182),
    .a({net_1038,net_247}),
    .b({net_1299,net_929}),
    .c({open_n553,net_1038}),
    .mi({open_n554,io_i2c_sda}),
    .f({net_826,net_825}),
    .q({open_n555,net_827})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hFF4F"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h5F00"),
    .INIT_LUTG1("16'h1300"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_441
  (
    .clk(gclk_9),
    .ce(net_454),
    .a({net_906,net_821}),
    .b({net_956,net_1283}),
    .c({net_946,net_312}),
    .d({net_822,net_1035}),
    .e({net_547,net_1286}),
    .mi({open_n556,io_mcu_d[0]}),
    .f({net_824,net_822}),
    .q({open_n557,net_821})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0A00"),
    .INIT_LUT1("16'hFF0B"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_442
  (
    .clk(gclk_9),
    .a({io_mcu_d[6],io_mcu_d[6]}),
    .b({net_265,net_793}),
    .c({i_mcu_dcs,i_mcu_dcs}),
    .d({net_793,net_265}),
    .mi({open_n558,net_823}),
    .q({open_n559,net_823})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h2222"),
    .INIT_LUTF1("16'hA888"),
    .INIT_LUTG1("16'hA888"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_443
  (
    .clk(gclk_8),
    .ce(net_830),
    .sr(net_182),
    .a({net_960,net_960}),
    .b({net_1303,net_247}),
    .c({net_962,open_n560}),
    .d({net_1289,open_n561}),
    .e({open_n562,net_1303}),
    .mi({open_n563,io_i2c_sda}),
    .f({net_829,net_830}),
    .q({open_n564,net_828})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h00A0"),
    .INIT_LUT1("16'h5F13"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_444
  (
    .clk(gclk_8),
    .ce(net_837),
    .sr(net_182),
    .a({net_1521,net_847}),
    .b({net_1525,open_n565}),
    .c({net_847,net_1521}),
    .d({net_952,net_247}),
    .mi({open_n566,io_i2c_sda}),
    .f({net_841,net_837}),
    .q({open_n567,net_833})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h2222"),
    .INIT_LUTF1("16'h5500"),
    .INIT_LUTG1("16'h0500"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_445
  (
    .clk(gclk_8),
    .ce(net_834),
    .sr(net_182),
    .a({net_684,net_1047}),
    .b({open_n568,net_247}),
    .c({net_1528,open_n569}),
    .d({net_846,open_n570}),
    .e({net_964,net_964}),
    .mi({open_n571,io_i2c_sda}),
    .f({net_836,net_834}),
    .q({open_n572,net_835})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h4444"),
    .INIT_LUTF1("16'h5500"),
    .INIT_LUTG1("16'h1100"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_446
  (
    .clk(gclk_8),
    .ce(net_842),
    .sr(net_182),
    .a({net_352,net_247}),
    .b({net_862,net_847}),
    .d({net_247,open_n573}),
    .e({net_1523,net_1523}),
    .mi({open_n574,io_i2c_sda}),
    .f({net_838,net_842}),
    .q({open_n575,net_831})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hF000"),
    .INIT_LUT1("16'hC000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_447
  (
    .clk(gclk_8),
    .ce(net_839),
    .sr(net_182),
    .b({net_1289,open_n576}),
    .c({net_952,net_960}),
    .d({net_960,net_920}),
    .mi({open_n577,io_i2c_sda}),
    .f({net_840,net_839}),
    .q({open_n578,net_832})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hC0C0"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h3F3F"),
    .INIT_LUTG1("16'h003F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_448
  (
    .clk(gclk_8),
    .ce(net_844),
    .sr(net_182),
    .b({net_1333,net_1056}),
    .c({net_843,net_1333}),
    .d({net_1648,open_n579}),
    .e({net_966,net_247}),
    .mi({open_n580,io_i2c_sda}),
    .f({net_846,net_844}),
    .q({open_n581,net_845})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h1000"),
    .INIT_LUT1("16'h1000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_449
  (
    .a({net_1532,net_1301}),
    .b({net_1299,net_1299}),
    .c({net_1301,net_1300}),
    .d({net_1300,net_1532}),
    .f({net_847,net_843})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h001F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_450
  (
    .a({net_1060,net_1060}),
    .b({net_584,net_584}),
    .c({net_1276,net_1276}),
    .d({net_1066,net_1066}),
    .mi({open_n582,net_1073}),
    .fx({open_n583,net_848})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hF000"),
    .INIT_LUTG0("16'hF000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h0808"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_451
  (
    .a({net_856,open_n584}),
    .b({net_480,open_n585}),
    .c({net_475,net_1182}),
    .d({open_n586,net_1312}),
    .e({net_1192,open_n587}),
    .f({net_850,net_849})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h6804"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_452
  (
    .a({net_1532,net_1532}),
    .b({net_1299,net_1301}),
    .c({net_1301,net_1300}),
    .d({net_1300,net_1299}),
    .mi({open_n588,net_1289}),
    .fx({open_n589,net_853})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h001F"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h003F"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_453
  (
    .a({open_n590,net_843}),
    .b({net_584,net_1078}),
    .c({net_1067,net_1060}),
    .d({net_568,net_954}),
    .e({net_954,net_1064}),
    .f({net_854,net_852})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hFF55"),
    .INIT_LUTG0("16'h0011"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hFEFE"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_454
  (
    .a({net_950,net_951}),
    .b({net_959,net_1301}),
    .c({net_962,open_n591}),
    .d({open_n592,net_1299}),
    .e({net_1060,net_1060}),
    .f({net_851,net_857})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h8000"),
    .INIT_LUT1("16'h0700"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_455
  (
    .a({net_564,net_564}),
    .b({net_959,net_1532}),
    .c({net_970,net_1300}),
    .d({net_1073,net_1299}),
    .f({net_856,net_855})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'hD700"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_456
  (
    .a({net_1057,net_1057}),
    .b({net_1532,net_1532}),
    .c({net_1301,net_1301}),
    .d({net_852,net_852}),
    .mi({open_n593,net_861}),
    .fx({open_n594,net_860})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0555"),
    .INIT_LUTG0("16'h0111"),
    .INIT_LUTF1("16'hD0D0"),
    .INIT_LUTG1("16'h1010"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_457
  (
    .a({net_1301,net_858}),
    .b({net_1300,net_961}),
    .c({net_584,net_592}),
    .d({open_n595,net_668}),
    .e({net_1299,net_1303}),
    .f({net_858,net_859})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h020A"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_458
  (
    .a({net_859,net_859}),
    .b({net_959,net_959}),
    .c({net_564,net_965}),
    .d({net_965,net_564}),
    .mi({open_n596,net_970}),
    .fx({open_n597,net_861})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hF0F0"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hF0F0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_459
  (
    .c({net_959,net_959}),
    .e({net_1301,net_1301}),
    .f({net_863,net_862})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hAAAA"),
    .INIT_LUT1("16'hEA2A"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_460
  (
    .clk(gclk_9),
    .ce(net_1107),
    .a({io_mcu_d[0],net_864}),
    .b({io_mcu_d[1],io_mcu_d[0]}),
    .c({io_mcu_d[2],io_mcu_d[2]}),
    .d({net_864,io_mcu_d[1]}),
    .mi({open_n598,net_641}),
    .q({open_n599,net_864})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h8AFA"),
    .INIT_LUT1("16'hA2EE"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_461
  (
    .clk(gclk_9),
    .ce(net_1107),
    .a({net_865,net_866}),
    .b({net_641,io_mcu_d[2]}),
    .c({io_mcu_d[1],net_641}),
    .d({io_mcu_d[2],io_mcu_d[1]}),
    .q({net_865,net_866})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h1155"),
    .INIT_LUTG0("16'h1100"),
    .INIT_LUTF1("16'h1155"),
    .INIT_LUTG1("16'h0044"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_466
  (
    .a({net_189,net_189}),
    .b({net_1044,net_701}),
    .d({net_699,net_1044}),
    .e({net_694,net_691}),
    .f({net_869,net_868})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h33AA"),
    .INIT_LUT1("16'h5555"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_467
  (
    .clk(gclk_4),
    .a({net_511,net_867}),
    .b({net_631,net_631}),
    .c({net_994,net_511}),
    .d({net_867,net_994}),
    .mi({open_n600,net_445}),
    .q({open_n601,net_867})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h33AA"),
    .INIT_LUT1("16'h0F0F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_468
  (
    .clk(gclk_4),
    .a({net_994,net_870}),
    .b({net_624,net_624}),
    .c({net_511,net_511}),
    .d({net_870,net_994}),
    .mi({open_n602,net_445}),
    .q({open_n603,net_870})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0545"),
    .INIT_LUTG0("16'h5545"),
    .INIT_LUTF1("16'h050F"),
    .INIT_LUTG1("16'h000A"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_469
  (
    .clk(gclk_4),
    .a({net_1044,net_871}),
    .b({open_n604,net_1537}),
    .c({net_189,net_189}),
    .d({net_703,net_1044}),
    .e({net_693,net_1546}),
    .mi({open_n605,net_1233}),
    .f({net_871,net_873}),
    .q({open_n606,net_872})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hAFCF"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_470
  (
    .a({net_1547,net_1547}),
    .b({net_1536,net_1536}),
    .c({net_189,net_189}),
    .d({net_1044,net_1044}),
    .mi({open_n607,net_219}),
    .fx({open_n608,net_874})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hCCAA"),
    .INIT_LUT1("16'h0F0F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_471
  (
    .clk(gclk_4),
    .a({net_994,net_875}),
    .b({net_876,net_876}),
    .c({net_511,net_511}),
    .d({net_875,net_994}),
    .mi({open_n609,net_445}),
    .q({open_n610,net_875})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h5555"),
    .INIT_LUTG0("16'hD555"),
    .INIT_LUTF1("16'h0001"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_472
  (
    .clk(gclk_5),
    .sr(net_880),
    .a({net_877,net_879}),
    .b({net_760,net_605}),
    .c({net_772,net_744}),
    .d({net_878,net_782}),
    .e({net_762,net_767}),
    .mi({net_766,net_769}),
    .f({net_879,net_880}),
    .q({net_877,net_878})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h33AA"),
    .INIT_LUT1("16'h3333"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_473
  (
    .clk(gclk_4),
    .a({net_623,net_876}),
    .b({net_511,net_623}),
    .c({net_994,net_511}),
    .d({net_876,net_994}),
    .mi({open_n611,net_445}),
    .q({open_n612,net_876})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h8000"),
    .INIT_LUT1("16'h0505"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_474
  (
    .clk(gclk_9),
    .ce(net_882),
    .a({net_881,net_222}),
    .b({open_n613,net_308}),
    .c({net_630,net_180}),
    .d({open_n614,net_181}),
    .mi({io_mcu_d[2],io_mcu_d[0]}),
    .f({net_883,net_882}),
    .q({net_881,net_884})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h00D0"),
    .INIT_LUTG0("16'hD0D0"),
    .INIT_LUTF1("16'h4400"),
    .INIT_LUTG1("16'h4F00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_475
  (
    .clk(gclk_9),
    .ce(net_779),
    .a({net_887,net_886}),
    .b({net_762,net_772}),
    .c({net_885,net_891}),
    .d({net_891,net_887}),
    .e({net_878,net_762}),
    .mi({io_mcu_d[4],io_mcu_d[7]}),
    .f({net_889,net_893}),
    .q({net_887,net_886})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hCF0C"),
    .INIT_LUTG0("16'hDF0D"),
    .INIT_LUTF1("16'h00F5"),
    .INIT_LUTG1("16'hF5F5"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_476
  (
    .clk(gclk_9),
    .ce(net_779),
    .a({net_885,net_888}),
    .b({open_n615,net_889}),
    .c({net_878,net_886}),
    .d({net_888,net_772}),
    .e({net_877,net_877}),
    .mi({io_mcu_d[5],io_mcu_d[6]}),
    .f({net_891,net_894}),
    .q({net_885,net_888})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h5555"),
    .INIT_LUT1("16'h007F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_477
  (
    .clk(gclk_5),
    .ce(net_785),
    .a({net_1353,net_890}),
    .b({net_1359,open_n616}),
    .c({net_1351,open_n617}),
    .d({net_1355,open_n618}),
    .f({net_892,open_n619}),
    .q({open_n620,net_890})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h1000"),
    .INIT_LUT1("16'hF000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_478
  (
    .clk(gclk_9),
    .ce(net_897),
    .a({open_n621,net_180}),
    .b({open_n622,net_181}),
    .c({net_533,net_1111}),
    .d({net_452,net_895}),
    .mi({io_mcu_d[3],io_mcu_d[0]}),
    .f({net_895,net_897}),
    .q({net_899,net_898})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h4000"),
    .INIT_LUTF1("16'h5050"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_479
  (
    .clk(gclk_9),
    .ce(net_900),
    .a({net_644,net_181}),
    .b({open_n623,net_1111}),
    .c({net_536,net_536}),
    .d({open_n624,net_180}),
    .e({net_643,net_452}),
    .mi({open_n625,io_mcu_d[0]}),
    .f({net_896,net_900}),
    .q({open_n626,net_901})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h2277"),
    .INIT_LUTG0("16'h2277"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h3F3F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_480
  (
    .a({open_n627,net_516}),
    .b({net_1341,net_987}),
    .c({net_908,open_n628}),
    .d({open_n629,net_179}),
    .e({net_1095,open_n630}),
    .f({net_902,net_903})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h8080"),
    .INIT_LUT1("16'h00C0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_481
  (
    .a({open_n631,net_180}),
    .b({net_181,net_181}),
    .c({net_896,net_896}),
    .d({net_180,open_n632}),
    .f({net_905,net_904})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h1000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_482
  (
    .a({net_180,net_180}),
    .b({net_181,net_181}),
    .c({net_647,net_647}),
    .d({net_644,net_644}),
    .mi({open_n633,net_643}),
    .fx({open_n634,net_906})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h4040"),
    .INIT_LUT1("16'h0777"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_483
  (
    .clk(gclk_8),
    .ce(net_912),
    .sr(net_182),
    .a({net_1209,net_247}),
    .b({net_905,net_943}),
    .c({net_648,net_1303}),
    .d({net_907,open_n635}),
    .mi({open_n636,io_i2c_sda}),
    .f({net_915,net_912}),
    .q({open_n637,net_907})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hCC55"),
    .INIT_LUTG0("16'hF0F0"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h4000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_484
  (
    .clk(gclk_9),
    .a({net_650,net_910}),
    .b({net_790,net_180}),
    .c({net_824,net_911}),
    .d({net_1008,i_mcu_dcs}),
    .e({net_1136,i_mcu_rws}),
    .f({net_910,open_n638}),
    .q({open_n639,net_911})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hCC0F"),
    .INIT_LUT1("16'hFF00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_485
  (
    .clk(gclk_9),
    .a({net_1022,net_908}),
    .b({net_644,net_644}),
    .c({i_mcu_dcs,net_1022}),
    .d({net_908,i_mcu_dcs}),
    .mi({open_n640,i_mcu_rws}),
    .q({open_n641,net_908})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h00AA"),
    .INIT_LUTF1("16'h0FFF"),
    .INIT_LUTG1("16'h0555"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_486
  (
    .clk(gclk_8),
    .ce(net_914),
    .sr(net_182),
    .a({net_1554,net_943}),
    .c({net_648,open_n642}),
    .d({net_909,net_247}),
    .e({net_904,net_1528}),
    .mi({open_n643,io_i2c_sda}),
    .f({net_913,net_914}),
    .q({open_n644,net_909})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h5000"),
    .INIT_LUT1("16'h4444"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_487
  (
    .clk(gclk_9),
    .ce(net_1149),
    .a({net_1283,net_1141}),
    .b({net_1349,open_n645}),
    .c({open_n646,net_911}),
    .d({open_n647,net_916}),
    .mi({open_n648,io_mcu_d[6]}),
    .f({net_916,net_918}),
    .q({open_n649,net_917})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hCCAA"),
    .INIT_LUTG0("16'hCCAA"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hFC0C"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_488
  (
    .clk(gclk_4),
    .ce(net_1291),
    .sr(net_445),
    .a({open_n650,net_1273}),
    .b({net_324,net_1176}),
    .c({net_1141,open_n651}),
    .d({net_919,net_527}),
    .e({net_439,open_n652}),
    .mi({open_n653,net_1273}),
    .f({net_922,net_921}),
    .q({open_n654,net_919})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hFA0A"),
    .INIT_LUT1("16'h11DD"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_489
  (
    .clk(gclk_4),
    .ce(net_1291),
    .sr(net_445),
    .a({net_736,net_1275}),
    .b({net_1044,open_n655}),
    .c({open_n656,net_527}),
    .d({net_727,net_1175}),
    .mi({open_n657,net_1275}),
    .f({net_925,net_924}),
    .q({open_n658,net_927})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h00A0"),
    .INIT_LUTG0("16'h00A0"),
    .INIT_LUTF1("16'h00AA"),
    .INIT_LUTG1("16'h00AA"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_490
  (
    .clk(gclk_8),
    .ce(net_926),
    .sr(net_182),
    .a({net_1528,net_1056}),
    .c({open_n659,net_1032}),
    .d({net_247,net_247}),
    .mi({open_n660,io_i2c_sda}),
    .f({net_920,net_926}),
    .q({open_n661,net_923})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hF0F0"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_491
  (
    .c({open_n662,net_963}),
    .f({open_n663,net_935})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0AAA"),
    .INIT_LUTG0("16'h0222"),
    .INIT_LUTF1("16'h7777"),
    .INIT_LUTG1("16'h0707"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_492
  (
    .clk(gclk_4),
    .a({net_832,net_930}),
    .b({net_796,i_adc1B_d[6]}),
    .c({net_999,net_1244}),
    .d({open_n664,i_adc1A_d[6]}),
    .e({net_833,net_794}),
    .mi({i_adc1A_d[6],i_adc1B_d[6]}),
    .f({net_930,net_931}),
    .q({net_933,net_938})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h3000"),
    .INIT_LUT1("16'h0004"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_493
  (
    .clk(gclk_8),
    .ce(net_934),
    .sr(net_182),
    .a({net_1532,open_n665}),
    .b({net_1299,net_247}),
    .c({net_1300,net_584}),
    .d({net_1301,net_929}),
    .mi({open_n666,io_i2c_sda}),
    .f({net_929,net_934}),
    .q({open_n667,net_932})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h1000"),
    .INIT_LUTF1("16'h33FF"),
    .INIT_LUTG1("16'h030F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_494
  (
    .clk(gclk_8),
    .ce(net_937),
    .sr(net_182),
    .a({open_n668,net_1302}),
    .b({net_998,net_247}),
    .c({net_999,net_1303}),
    .d({net_928,net_948}),
    .e({net_676,net_963}),
    .mi({open_n669,io_i2c_sda}),
    .f({net_936,net_937}),
    .q({open_n670,net_928})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0A00"),
    .INIT_LUT1("16'hAA00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_495
  (
    .clk(gclk_8),
    .ce(net_940),
    .sr(net_182),
    .a({net_1067,net_584}),
    .c({open_n671,net_247}),
    .d({net_1289,net_1067}),
    .mi({open_n672,io_i2c_sda}),
    .f({net_939,net_940}),
    .q({open_n673,net_941})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0777"),
    .INIT_LUTF1("16'hFF00"),
    .INIT_LUTG1("16'h5500"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_496
  (
    .clk(gclk_4),
    .a({net_906,net_794}),
    .b({open_n674,i_adc1B_d[1]}),
    .c({open_n675,net_547}),
    .d({net_942,net_835}),
    .e({net_577,net_1013}),
    .mi({open_n676,i_adc1B_d[1]}),
    .f({net_947,net_942}),
    .q({open_n677,net_944})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'hAAAA"),
    .INIT_LUTF1("16'h0030"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_497
  (
    .clk(gclk_8),
    .ce(net_945),
    .sr(net_182),
    .a({open_n678,net_920}),
    .b({net_948,open_n679}),
    .c({net_1182,open_n680}),
    .d({net_1312,open_n681}),
    .e({net_1302,net_1525}),
    .mi({open_n682,io_i2c_sda}),
    .f({net_943,net_945}),
    .q({open_n683,net_946})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h4000"),
    .INIT_LUT1("16'hF000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_498
  (
    .clk(gclk_8),
    .ce(net_1530),
    .sr(net_182),
    .a({open_n684,net_948}),
    .b({open_n685,net_963}),
    .c({net_1329,net_1302}),
    .d({net_939,net_939}),
    .mi({open_n686,net_1310}),
    .f({net_957,net_954}),
    .q({open_n687,net_948})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h00AA"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hAAAA"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_499
  (
    .clk(gclk_8),
    .ce(net_953),
    .sr(net_182),
    .a({net_964,net_964}),
    .d({open_n688,net_247}),
    .e({net_1289,net_1303}),
    .mi({open_n689,io_i2c_sda}),
    .f({net_951,net_953}),
    .q({open_n690,net_956})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0003"),
    .INIT_LUTG0("16'h00FF"),
    .INIT_LUTF1("16'hA0A0"),
    .INIT_LUTG1("16'hF0F0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_500
  (
    .a({net_939,open_n691}),
    .b({open_n692,net_1303}),
    .c({net_1648,net_1528}),
    .d({open_n693,net_949}),
    .e({net_1528,net_1159}),
    .f({net_949,net_955})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h8000"),
    .INIT_LUT1("16'h4000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_501
  (
    .a({net_1299,net_1532}),
    .b({net_1532,net_1301}),
    .c({net_1300,net_1300}),
    .d({net_1301,net_1299}),
    .f({net_950,net_952})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h001F"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_502
  (
    .a({net_950,net_950}),
    .b({net_668,net_847}),
    .c({net_847,net_668}),
    .d({net_855,net_855}),
    .mi({open_n694,net_1500}),
    .fx({open_n695,net_958})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h00AA"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h5500"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_503
  (
    .a({net_948,net_948}),
    .d({net_1302,net_1302}),
    .e({net_849,net_849}),
    .f({net_960,net_961})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h2000"),
    .INIT_LUTG0("16'h2000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h2222"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_504
  (
    .a({net_1532,net_1299}),
    .b({net_1300,net_1301}),
    .c({open_n696,net_1532}),
    .d({open_n697,net_1300}),
    .e({net_1299,open_n698}),
    .f({net_959,net_962})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hA000"),
    .INIT_LUT1("16'hA0A0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_505
  (
    .a({net_470,net_1329}),
    .c({net_1329,net_1289}),
    .d({open_n699,net_592}),
    .f({net_965,net_969})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0055"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h8888"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_506
  (
    .a({net_1302,net_948}),
    .b({net_948,open_n700}),
    .d({open_n701,net_1302}),
    .e({net_849,net_849}),
    .f({net_967,net_964})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hAA00"),
    .INIT_LUTG0("16'hAA00"),
    .INIT_LUTF1("16'h0033"),
    .INIT_LUTG1("16'h0033"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_507
  (
    .a({open_n702,net_1289}),
    .b({net_1182,open_n703}),
    .d({net_1312,net_585}),
    .f({net_963,net_966})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h4000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_508
  (
    .a({net_948,net_948}),
    .b({net_963,net_963}),
    .c({net_1289,net_1289}),
    .d({net_1302,net_1302}),
    .mi({open_n704,net_592}),
    .fx({open_n705,net_968})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h1337"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_509
  (
    .a({net_1532,net_1532}),
    .b({net_1299,net_1301}),
    .c({net_1301,net_1300}),
    .d({net_1300,net_1299}),
    .mi({open_n706,net_1523}),
    .fx({open_n707,net_970})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hAAAA"),
    .INIT_LUT1("16'hEA2A"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_510
  (
    .clk(gclk_9),
    .ce(net_1117),
    .a({io_mcu_d[0],net_971}),
    .b({io_mcu_d[1],io_mcu_d[0]}),
    .c({io_mcu_d[2],io_mcu_d[2]}),
    .d({net_971,io_mcu_d[1]}),
    .mi({open_n708,net_641}),
    .q({open_n709,net_971})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hFAFA"),
    .INIT_LUTG0("16'h8A8A"),
    .INIT_LUTF1("16'hFAFA"),
    .INIT_LUTG1("16'h8A8A"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_511
  (
    .clk(gclk_9),
    .ce(net_1117),
    .a({net_973,net_972}),
    .b({io_mcu_d[1],io_mcu_d[2]}),
    .c({net_641,net_641}),
    .e({io_mcu_d[2],io_mcu_d[1]}),
    .q({net_973,net_972})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hCCAA"),
    .INIT_LUT1("16'h3333"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_512
  (
    .clk(gclk_4),
    .a({net_867,net_974}),
    .b({net_511,net_867}),
    .c({net_994,net_511}),
    .d({net_974,net_994}),
    .mi({open_n710,net_445}),
    .q({open_n711,net_974})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hFCFF"),
    .INIT_LUTG0("16'hC0CC"),
    .INIT_LUTF1("16'hAA00"),
    .INIT_LUTG1("16'hAA00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_513
  (
    .a({net_881,open_n712}),
    .b({open_n713,net_746}),
    .c({open_n714,net_982}),
    .d({net_630,net_884}),
    .e({open_n715,net_978}),
    .f({net_975,net_976})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h5440"),
    .INIT_LUT1("16'h5454"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_514
  (
    .a({net_1097,net_1097}),
    .b({net_631,net_631}),
    .c({net_1085,net_1085}),
    .d({net_975,net_975}),
    .mi({open_n716,net_980}),
    .fx({open_n717,net_977})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0077"),
    .INIT_LUTG0("16'h0017"),
    .INIT_LUTF1("16'h0E08"),
    .INIT_LUTG1("16'h0F0C"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_515
  (
    .clk(gclk_9),
    .ce(net_882),
    .a({net_781,net_978}),
    .b({net_636,net_636}),
    .c({net_883,net_781}),
    .d({net_978,net_975}),
    .e({net_884,net_884}),
    .mi({open_n718,io_mcu_d[1]}),
    .f({net_980,net_979}),
    .q({open_n719,net_978})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h33AA"),
    .INIT_LUT1("16'h0F0F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_516
  (
    .clk(gclk_4),
    .a({net_994,net_981}),
    .b({net_630,net_630}),
    .c({net_511,net_511}),
    .d({net_981,net_994}),
    .mi({open_n720,net_445}),
    .q({open_n721,net_981})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0545"),
    .INIT_LUTG0("16'h5545"),
    .INIT_LUTF1("16'h00AF"),
    .INIT_LUTG1("16'h0005"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_517
  (
    .clk(gclk_4),
    .a({net_1044,net_984}),
    .b({open_n722,net_1541}),
    .c({net_695,net_189}),
    .d({net_189,net_1044}),
    .e({net_707,net_1551}),
    .mi({open_n723,net_1232}),
    .f({net_984,net_987}),
    .q({open_n724,net_988})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h003F"),
    .INIT_LUTG0("16'h005F"),
    .INIT_LUTF1("16'h3000"),
    .INIT_LUTG1("16'h3033"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_518
  (
    .clk(gclk_4),
    .a({open_n725,net_1550}),
    .b({net_189,net_1542}),
    .c({net_706,net_189}),
    .d({net_1044,net_983}),
    .e({net_696,net_1044}),
    .mi({open_n726,net_1223}),
    .f({net_983,net_985}),
    .q({open_n727,net_986})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hCCAA"),
    .INIT_LUT1("16'h3333"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_519
  (
    .clk(gclk_4),
    .a({net_989,net_982}),
    .b({net_511,net_989}),
    .c({net_994,net_511}),
    .d({net_982,net_994}),
    .mi({open_n728,net_445}),
    .q({open_n729,net_982})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hF4FF"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("INV"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_520
  (
    .clk(gclk_5),
    .ce(net_880),
    .a({open_n730,net_760}),
    .b({open_n731,net_776}),
    .c({open_n732,net_784}),
    .d({open_n733,net_893}),
    .e({open_n734,net_894}),
    .q({open_n735,net_990})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h33AA"),
    .INIT_LUT1("16'h5555"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_521
  (
    .clk(gclk_4),
    .a({net_511,net_989}),
    .b({net_781,net_781}),
    .c({net_994,net_511}),
    .d({net_989,net_994}),
    .mi({open_n736,net_445}),
    .q({open_n737,net_989})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h5F3F"),
    .INIT_LUTF1("16'hCE0E"),
    .INIT_LUTG1("16'hEEAE"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_522
  (
    .clk(gclk_4),
    .a({net_991,net_1549}),
    .b({net_614,net_1540}),
    .c({net_523,net_904}),
    .d({net_1048,net_1044}),
    .e({net_629,net_189}),
    .mi({open_n738,net_1226}),
    .f({net_993,net_991}),
    .q({open_n739,net_992})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h000A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD_CARRY"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("F"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_523
  (
    .clk(gclk_5),
    .sr(net_785),
    .a({net_996,1'b0}),
    .q({net_996,open_n740}),
    .fco(block_523_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_525
  (
    .clk(gclk_5),
    .sr(net_785),
    .a({net_995,net_997}),
    .b({1'b0,1'b0}),
    .fci(block_523_carry),
    .q({net_995,net_997}),
    .fco(block_525_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_527
  (
    .clk(gclk_5),
    .sr(net_785),
    .a({net_1002,net_1005}),
    .b({1'b0,1'b0}),
    .fci(block_525_carry),
    .q({net_1002,net_1005}),
    .fco(block_527_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_529
  (
    .clk(gclk_5),
    .sr(net_785),
    .a({net_1001,net_1003}),
    .b({1'b0,1'b0}),
    .fci(block_527_carry),
    .q({net_1001,net_1003}),
    .fco(block_529_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_530
  (
    .clk(gclk_5),
    .sr(net_785),
    .a({open_n741,net_1009}),
    .b({open_n742,1'b0}),
    .fci(block_529_carry),
    .q({open_n743,net_1009})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hEEEE"),
    .INIT_LUTG0("16'hFFFF"),
    .INIT_LUTF1("16'hBBBB"),
    .INIT_LUTG1("16'h1111"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_524
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1044,net_994}),
    .b({net_710,net_1222}),
    .e({net_718,net_1241}),
    .f({net_1000,open_n744}),
    .q({open_n745,net_994})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h1010"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h4040"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_526
  (
    .a({net_180,net_180}),
    .b({net_181,net_181}),
    .c({net_647,net_647}),
    .e({net_1111,net_1111}),
    .f({net_999,net_998})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h1000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h002A"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_528
  (
    .clk(gclk_4),
    .a({net_780,net_1496}),
    .b({net_1167,net_180}),
    .c({net_796,net_309}),
    .d({net_1004,net_1111}),
    .e({net_1258,net_181}),
    .mi({i_adc1B_d[0],net_1227}),
    .f({net_1008,net_1004}),
    .q({net_1007,net_1006})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0007"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h5F5F"),
    .INIT_LUTG1("16'h005F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_531
  (
    .clk(gclk_4),
    .a({i_adc1A_d[1],net_1111}),
    .b({open_n746,net_647}),
    .c({net_1244,net_1244}),
    .d({i_adc2B_d[1],net_896}),
    .e({net_1242,net_796}),
    .mi({i_adc1A_d[1],i_adc2B_d[1]}),
    .f({net_1013,net_1010}),
    .q({net_1011,net_1012})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0088"),
    .INIT_LUT1("16'h153F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_532
  (
    .clk(gclk_8),
    .ce(net_1020),
    .sr(net_182),
    .a({net_998,net_1523}),
    .b({net_999,net_1067}),
    .c({net_1519,open_n747}),
    .d({net_1014,net_247}),
    .mi({open_n748,io_i2c_sda}),
    .f({net_1021,net_1020}),
    .q({open_n749,net_1014})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h4040"),
    .INIT_LUTG0("16'h4040"),
    .INIT_LUTF1("16'h55FF"),
    .INIT_LUTG1("16'h050F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_533
  (
    .clk(gclk_8),
    .ce(net_1018),
    .sr(net_182),
    .a({net_796,net_247}),
    .b({open_n750,net_847}),
    .c({net_999,net_584}),
    .d({net_1015,open_n751}),
    .e({net_1166,open_n752}),
    .mi({open_n753,io_i2c_sda}),
    .f({net_1017,net_1018}),
    .q({open_n754,net_1015})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0FBF"),
    .INIT_LUTF1("16'h8000"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_534
  (
    .clk(gclk_9),
    .ce(net_1156),
    .a({net_1016,net_1141}),
    .b({net_902,net_908}),
    .c({net_551,net_1349}),
    .d({net_815,net_1283}),
    .e({net_1028,net_1247}),
    .mi({open_n755,io_mcu_d[6]}),
    .f({net_1022,net_1016}),
    .q({open_n756,net_1019})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h00B0"),
    .INIT_LUT1("16'h0407"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_535
  (
    .clk(gclk_4),
    .ce(net_1291),
    .sr(net_445),
    .a({net_1152,net_1025}),
    .b({net_1141,net_1283}),
    .c({net_1283,net_439}),
    .d({net_908,net_1023}),
    .mi({open_n757,net_1279}),
    .f({net_1023,net_1028}),
    .q({open_n758,net_1025})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0808"),
    .INIT_LUTG0("16'h0808"),
    .INIT_LUTF1("16'h33FF"),
    .INIT_LUTG1("16'h030F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_536
  (
    .clk(gclk_8),
    .ce(net_1027),
    .sr(net_182),
    .a({open_n759,net_1067}),
    .b({net_547,net_951}),
    .c({net_923,net_247}),
    .d({net_1024,open_n760}),
    .e({net_906,open_n761}),
    .mi({open_n762,io_i2c_sda}),
    .f({net_1026,net_1027}),
    .q({open_n763,net_1024})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hE0E0"),
    .INIT_LUTG0("16'hEEAA"),
    .INIT_LUTF1("16'hF0CC"),
    .INIT_LUTG1("16'hF0CC"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_537
  (
    .clk(gclk_4),
    .ce(net_1291),
    .sr(net_445),
    .a({open_n764,net_916}),
    .b({net_1274,net_439}),
    .c({net_1181,net_256}),
    .d({net_527,net_1029}),
    .e({open_n765,net_1141}),
    .mi({net_1274,open_n766}),
    .f({net_1031,net_1030}),
    .q({net_1029,open_n767})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h2200"),
    .INIT_LUT1("16'hA0A0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_538
  (
    .clk(gclk_8),
    .ce(net_1040),
    .sr(net_182),
    .a({net_1289,net_1276}),
    .b({open_n768,net_247}),
    .c({net_1525,open_n769}),
    .d({open_n770,net_1032}),
    .mi({open_n771,io_i2c_sda}),
    .f({net_1032,net_1040}),
    .q({open_n772,net_1043})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h4040"),
    .INIT_LUTF1("16'hA000"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_539
  (
    .clk(gclk_8),
    .ce(net_1036),
    .sr(net_182),
    .a({net_935,net_1302}),
    .b({open_n773,net_963}),
    .c({net_1289,net_948}),
    .d({net_948,open_n774}),
    .e({net_1302,net_920}),
    .mi({open_n775,io_i2c_sda}),
    .f({net_1038,net_1036}),
    .q({open_n776,net_1042})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h050F"),
    .INIT_LUTG0("16'h0500"),
    .INIT_LUTF1("16'hAA88"),
    .INIT_LUTG1("16'h2200"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_540
  (
    .a({net_896,net_1180}),
    .b({net_180,open_n777}),
    .c({open_n778,i_mcu_rws}),
    .d({net_95,net_896}),
    .e({net_329,net_1330}),
    .f({net_1041,net_1033})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0503"),
    .INIT_LUT1("16'h0407"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_541
  (
    .clk(gclk_9),
    .ce(net_1149),
    .a({net_538,net_1297}),
    .b({net_1141,net_911}),
    .c({net_1283,net_1283}),
    .d({net_911,net_1141}),
    .mi({io_mcu_d[5],io_mcu_d[2]}),
    .f({net_1035,net_1034}),
    .q({net_1037,net_1039})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h000A"),
    .INIT_LUTG0("16'h0002"),
    .INIT_LUTF1("16'h33FF"),
    .INIT_LUTG1("16'h1155"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_542
  (
    .clk(gclk_4),
    .a({i_adc1A_d[4],net_1045}),
    .b({net_1058,i_adc1B_d[4]}),
    .c({open_n779,net_922}),
    .d({net_796,net_241}),
    .e({net_1244,net_794}),
    .mi({i_adc1A_d[4],i_adc1B_d[4]}),
    .f({net_1045,net_1049}),
    .q({net_1046,net_1051})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hEE44"),
    .INIT_LUT1("16'h5533"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_543
  (
    .clk(gclk_3),
    .a({net_726,net_527}),
    .b({net_735,net_1279}),
    .d({net_1044,net_1195}),
    .f({net_1048,net_1050}),
    .q({open_n780,net_1044})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h0040"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_544
  (
    .a({net_1532,net_1532}),
    .b({net_1289,net_1300}),
    .c({net_1301,net_1301}),
    .d({net_1300,net_1289}),
    .mi({open_n781,net_1299}),
    .fx({open_n782,net_1047})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h8888"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h8080"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_545
  (
    .clk(gclk_8),
    .ce(net_1054),
    .sr(net_182),
    .a({net_1314,net_929}),
    .b({net_1287,net_1032}),
    .c({net_1186,open_n783}),
    .e({net_1055,net_247}),
    .mi({open_n784,io_i2c_sda}),
    .f({net_1052,net_1054}),
    .q({open_n785,net_1053})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hFFFF"),
    .INIT_LUT1("16'hFF70"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_546
  (
    .clk(gclk_8),
    .sr(net_182),
    .a({net_247,net_247}),
    .b({net_1055,net_1055}),
    .c({net_1186,net_1186}),
    .d({net_1189,net_1189}),
    .mi({open_n786,net_1295}),
    .q({open_n787,net_1062})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h8888"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h0C0C"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_547
  (
    .clk(gclk_8),
    .ce(net_1061),
    .sr(net_182),
    .a({open_n788,net_1056}),
    .b({net_1301,net_584}),
    .c({net_1532,open_n789}),
    .e({net_1077,net_247}),
    .mi({open_n790,io_i2c_sda}),
    .f({net_1056,net_1061}),
    .q({open_n791,net_1058})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h8888"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hCCCC"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_548
  (
    .clk(gclk_8),
    .ce(net_1063),
    .sr(net_182),
    .a({open_n792,net_1333}),
    .b({net_1333,net_1067}),
    .e({net_1077,net_247}),
    .mi({open_n793,io_i2c_sda}),
    .f({net_1057,net_1063}),
    .q({open_n794,net_1059})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0044"),
    .INIT_LUT1("16'hAA00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_549
  (
    .a({net_1055,net_948}),
    .b({open_n795,net_963}),
    .d({net_1289,net_1302}),
    .f({net_1060,net_1055})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hAA33"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h00AA"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_550
  (
    .a({net_963,net_1057}),
    .b({open_n796,net_1055}),
    .d({net_948,net_1532}),
    .e({net_966,net_966}),
    .f({net_1064,net_1065})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'hF888"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_551
  (
    .a({net_1303,net_1303}),
    .b({net_961,net_961}),
    .c({net_670,net_670}),
    .d({net_967,net_967}),
    .mi({open_n797,net_247}),
    .fx({open_n798,net_1066})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0A0A"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h8888"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_552
  (
    .a({net_1077,net_1077}),
    .b({net_584,open_n799}),
    .c({open_n800,net_1301}),
    .e({net_1301,net_1532}),
    .f({net_1068,net_1067})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0545"),
    .INIT_LUTG0("16'h5545"),
    .INIT_LUTF1("16'h4477"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("INV"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_553
  (
    .clk(gclk_9),
    .ce(i_mcu_dcs),
    .a({net_1191,net_1072}),
    .b({net_896,net_1070}),
    .c({open_n801,i_mcu_rws}),
    .d({net_1070,net_453}),
    .e({i_mcu_rws,io_mcu_d[2]}),
    .f({net_1072,open_n802}),
    .q({open_n803,net_1070})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h00AF"),
    .INIT_LUTG0("16'h00CF"),
    .INIT_LUTF1("16'h0A0F"),
    .INIT_LUTG1("16'h0005"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("INV"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_554
  (
    .clk(gclk_9),
    .ce(i_mcu_dcs),
    .a({net_896,net_1069}),
    .b({open_n804,io_mcu_d[0]}),
    .c({i_mcu_rws,i_mcu_rws}),
    .d({net_1069,net_1071}),
    .e({net_1194,net_453}),
    .f({net_1071,open_n805}),
    .q({open_n806,net_1069})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h7F7F"),
    .INIT_LUT1("16'h070F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_555
  (
    .a({net_963,net_1302}),
    .b({net_470,net_470}),
    .c({net_1521,net_963}),
    .d({net_1302,net_1521}),
    .mi({open_n807,net_847}),
    .fx({open_n808,net_1073})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0055"),
    .INIT_LUT1("16'hA0A0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_556
  (
    .a({net_1077,net_1299}),
    .c({net_1532,open_n809}),
    .d({open_n810,net_1300}),
    .f({net_1078,net_1077})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0545"),
    .INIT_LUTG0("16'h5545"),
    .INIT_LUTF1("16'h0A0F"),
    .INIT_LUTG1("16'h0005"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("INV"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_557
  (
    .clk(gclk_9),
    .ce(i_mcu_dcs),
    .a({net_896,net_1076}),
    .b({open_n811,net_1075}),
    .c({i_mcu_rws,i_mcu_rws}),
    .d({net_1075,net_453}),
    .e({net_1188,io_mcu_d[1]}),
    .f({net_1076,open_n812}),
    .q({open_n813,net_1075})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hCFAF"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("INV"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_558
  (
    .clk(gclk_9),
    .ce(i_mcu_dcs),
    .a({net_453,net_1074}),
    .b({io_mcu_d[3],io_mcu_d[3]}),
    .c({i_mcu_rws,i_mcu_rws}),
    .d({net_1074,net_453}),
    .mi({open_n814,net_1201}),
    .q({open_n815,net_1074})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hBBB0"),
    .INIT_LUT1("16'hB000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_559
  (
    .a({net_974,net_974}),
    .b({net_1085,net_1085}),
    .c({net_976,net_976}),
    .d({net_1205,net_1205}),
    .mi({open_n816,net_881}),
    .fx({open_n817,net_1081})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hF351"),
    .INIT_LUTG0("16'h5100"),
    .INIT_LUTF1("16'hF0F0"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_560
  (
    .a({open_n818,net_1080}),
    .b({open_n819,net_1205}),
    .c({net_982,net_881}),
    .d({open_n820,net_978}),
    .e({net_884,net_746}),
    .f({net_1080,net_1082})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hCCAA"),
    .INIT_LUT1("16'h3333"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_561
  (
    .clk(gclk_4),
    .a({net_870,net_1079}),
    .b({net_511,net_870}),
    .c({net_994,net_511}),
    .d({net_1079,net_994}),
    .mi({open_n821,net_445}),
    .q({open_n822,net_1079})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hAFCF"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_562
  (
    .a({net_1543,net_1543}),
    .b({net_1535,net_1535}),
    .c({net_1044,net_189}),
    .d({net_189,net_1044}),
    .mi({open_n823,net_868}),
    .fx({open_n824,net_1083})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h7771"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0701"),
    .INIT_LUTG1("16'h0707"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_563
  (
    .clk(gclk_9),
    .ce(net_882),
    .a({net_1086,net_1085}),
    .b({net_624,net_631}),
    .c({net_1098,net_979}),
    .d({net_1087,net_883}),
    .e({net_1097,net_1099}),
    .mi({io_mcu_d[5],io_mcu_d[3]}),
    .f({net_1089,net_1087}),
    .q({net_1086,net_1085})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h00E8"),
    .INIT_LUTG0("16'h00FC"),
    .INIT_LUTF1("16'h00FF"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_564
  (
    .a({open_n825,net_1099}),
    .b({open_n826,net_1086}),
    .c({open_n827,net_624}),
    .d({net_903,net_1088}),
    .e({net_1092,net_977}),
    .f({net_1088,net_1090})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h33AA"),
    .INIT_LUT1("16'h3333"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_565
  (
    .clk(gclk_4),
    .a({net_783,net_1084}),
    .b({net_511,net_783}),
    .c({net_994,net_511}),
    .d({net_1084,net_994}),
    .mi({open_n828,net_445}),
    .q({open_n829,net_1084})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0505"),
    .INIT_LUT1("16'hF000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_566
  (
    .clk(gclk_9),
    .ce(net_882),
    .a({open_n830,net_1091}),
    .c({net_783,net_783}),
    .d({net_1091,open_n831}),
    .mi({open_n832,io_mcu_d[4]}),
    .f({net_1099,net_1097}),
    .q({open_n833,net_1091})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h5F3F"),
    .INIT_LUTF1("16'hCE0E"),
    .INIT_LUTG1("16'hEEAE"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_567
  (
    .clk(gclk_4),
    .a({net_1093,net_1544}),
    .b({net_750,net_1534}),
    .c({net_523,net_904}),
    .d({net_925,net_1044}),
    .e({net_1000,net_189}),
    .mi({open_n834,net_1224}),
    .f({net_1095,net_1093}),
    .q({open_n835,net_1096})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h8888"),
    .INIT_LUT1("16'h8421"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_568
  (
    .clk(gclk_9),
    .ce(net_882),
    .a({net_875,net_1092}),
    .b({net_1482,net_903}),
    .c({net_1213,open_n836}),
    .d({net_1092,open_n837}),
    .mi({open_n838,io_mcu_d[6]}),
    .f({net_1094,net_1098}),
    .q({open_n839,net_1092})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h33AA"),
    .INIT_LUT1("16'h0F0F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_569
  (
    .clk(gclk_4),
    .a({net_903,net_1100}),
    .b({net_994,net_903}),
    .c({net_511,net_511}),
    .d({net_1100,net_994}),
    .mi({open_n840,net_445}),
    .q({open_n841,net_1100})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0005"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0CCC"),
    .INIT_LUTG1("16'h0CCC"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_570
  (
    .clk(gclk_4),
    .a({open_n842,net_1224}),
    .b({net_820,open_n843}),
    .c({net_794,net_1227}),
    .d({i_adc1B_d[7],net_1226}),
    .e({open_n844,net_1214}),
    .mi({i_adc1B_d[7],net_1214}),
    .f({net_1108,net_1105}),
    .q({net_1104,net_1103})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h1000"),
    .INIT_LUTF1("16'h00D4"),
    .INIT_LUTG1("16'hD4FF"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_571
  (
    .clk(gclk_9),
    .ce(net_897),
    .a({net_1101,net_644}),
    .b({net_1355,net_643}),
    .c({net_1229,net_181}),
    .d({net_1102,net_895}),
    .e({net_1358,net_180}),
    .mi({io_mcu_d[4],io_mcu_d[5]}),
    .f({net_1106,net_1107}),
    .q({net_1101,net_1102})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h0777"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_572
  (
    .a({net_905,net_905}),
    .b({net_1212,net_1212}),
    .c({net_904,net_904}),
    .d({net_1552,net_1552}),
    .mi({open_n845,net_1490}),
    .fx({open_n846,net_1114})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hDCFD"),
    .INIT_LUTG0("16'h40C4"),
    .INIT_LUTF1("16'h4400"),
    .INIT_LUTG1("16'hFFFF"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("INV"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_573
  (
    .clk(gclk_6),
    .ce(net_1112),
    .a({net_892,net_1106}),
    .b({net_1358,net_1109}),
    .c({open_n847,net_1110}),
    .d({net_1354,net_1354}),
    .e({net_1370,net_1370}),
    .f({net_1112,open_n848}),
    .q({open_n849,net_1118})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h3333"),
    .INIT_LUTF1("16'hF000"),
    .INIT_LUTG1("16'hF000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_574
  (
    .clk(gclk_9),
    .ce(net_897),
    .b({open_n850,net_644}),
    .c({net_895,open_n851}),
    .d({net_249,open_n852}),
    .e({open_n853,net_643}),
    .mi({io_mcu_d[6],io_mcu_d[7]}),
    .f({net_1117,net_1111}),
    .q({net_1110,net_1109})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h4000"),
    .INIT_LUT1("16'h8000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_575
  (
    .clk(gclk_9),
    .ce(net_1116),
    .a({net_180,net_180}),
    .b({net_647,net_222}),
    .c({net_1111,net_1111}),
    .d({net_181,net_181}),
    .mi({open_n854,io_mcu_d[0]}),
    .f({net_1113,net_1116}),
    .q({open_n855,net_1115})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0088"),
    .INIT_LUT1("16'h0777"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_576
  (
    .clk(gclk_8),
    .ce(net_1120),
    .sr(net_182),
    .a({net_904,net_929}),
    .b({net_1553,net_668}),
    .c({net_1113,open_n856}),
    .d({net_1119,net_247}),
    .mi({open_n857,io_i2c_sda}),
    .f({net_1121,net_1120}),
    .q({open_n858,net_1119})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h000A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD_CARRY"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_577
  (
    .clk(gclk_9),
    .ce(net_640),
    .a({net_1507,1'b0}),
    .mi({open_n859,io_mcu_d[0]}),
    .f({net_1129,open_n860}),
    .q({open_n861,net_1130}),
    .fco(block_577_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_579
  (
    .clk(gclk_9),
    .ce(net_1259),
    .a({net_1264,net_1263}),
    .b({1'b0,1'b0}),
    .mi({io_mcu_d[2],io_mcu_d[1]}),
    .fci(block_577_carry),
    .f({net_1127,net_1128}),
    .q({net_1124,net_1123}),
    .fco(block_579_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_580
  (
    .clk(gclk_9),
    .ce(net_1259),
    .a({open_n862,net_1508}),
    .b({open_n863,1'b0}),
    .mi({io_mcu_d[7],io_mcu_d[6]}),
    .fci(block_579_carry),
    .f({open_n864,net_1132}),
    .q({net_1137,net_1138})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h2020"),
    .INIT_LUTG0("16'h2020"),
    .INIT_LUTF1("16'hAA00"),
    .INIT_LUTG1("16'hAA00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_578
  (
    .clk(gclk_8),
    .ce(net_1126),
    .sr(net_182),
    .a({net_998,net_1056}),
    .b({open_n865,net_247}),
    .c({open_n866,net_1523}),
    .d({net_1122,open_n867}),
    .mi({open_n868,io_i2c_sda}),
    .f({net_1125,net_1126}),
    .q({open_n869,net_1122})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0AAA"),
    .INIT_LUTG0("16'h0222"),
    .INIT_LUTF1("16'h55FF"),
    .INIT_LUTG1("16'h050F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_581
  (
    .clk(gclk_4),
    .a({net_845,net_1131}),
    .b({open_n870,i_adc1A_d[0]}),
    .c({net_998,i_adc2B_d[0]}),
    .d({net_999,net_1242}),
    .e({net_831,net_1244}),
    .mi({open_n871,i_adc1A_d[0]}),
    .f({net_1131,net_1136}),
    .q({open_n872,net_1139})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h00F0"),
    .INIT_LUT1("16'h135F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_582
  (
    .clk(gclk_4),
    .a({i_adc1A_d[3],open_n873}),
    .b({i_adc1B_d[3],open_n874}),
    .c({net_1244,net_994}),
    .d({net_794,net_1348}),
    .mi({i_adc1B_d[3],net_1241}),
    .f({net_1135,net_1140}),
    .q({net_1134,net_1133})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0100"),
    .INIT_LUT1("16'hAA00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_583
  (
    .clk(gclk_9),
    .ce(net_1269),
    .a({net_1141,net_1263}),
    .b({open_n875,net_1264}),
    .c({open_n876,net_1508}),
    .d({net_525,net_1507}),
    .mi({open_n877,io_mcu_d[6]}),
    .f({net_1142,net_1141}),
    .q({open_n878,net_1143})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h4000"),
    .INIT_LUTF1("16'hCC00"),
    .INIT_LUTG1("16'hCC00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_584
  (
    .clk(gclk_9),
    .ce(net_1149),
    .a({open_n879,net_180}),
    .b({net_1141,net_224}),
    .c({open_n880,net_181}),
    .d({net_1145,net_644}),
    .e({open_n881,net_643}),
    .mi({io_mcu_d[0],io_mcu_d[1]}),
    .f({net_1149,net_1145}),
    .q({net_1151,net_1153})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hAA00"),
    .INIT_LUTG0("16'hAAFF"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hFA0A"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_585
  (
    .clk(gclk_4),
    .ce(net_1291),
    .sr(net_445),
    .a({net_190,net_1177}),
    .c({net_1141,open_n882}),
    .d({net_1144,net_527}),
    .e({net_439,net_1272}),
    .mi({open_n883,net_1272}),
    .f({net_1148,net_1147}),
    .q({open_n884,net_1144})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hFA0A"),
    .INIT_LUT1("16'hFA0A"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_586
  (
    .clk(gclk_4),
    .ce(net_1291),
    .sr(net_445),
    .a({net_1265,net_1282}),
    .c({net_527,net_527}),
    .d({net_1170,net_1187}),
    .mi({net_1265,net_1282}),
    .f({net_1146,net_1154}),
    .q({net_1152,net_1150})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hAACC"),
    .INIT_LUTG0("16'hF0F0"),
    .INIT_LUTF1("16'hC0C0"),
    .INIT_LUTG1("16'hC0C0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_587
  (
    .clk(gclk_9),
    .ce(net_1156),
    .a({open_n885,net_1293}),
    .b({net_1145,net_662}),
    .c({net_1283,net_1296}),
    .d({open_n886,net_1141}),
    .e({open_n887,net_1283}),
    .mi({io_mcu_d[0],io_mcu_d[5]}),
    .f({net_1156,net_1160}),
    .q({net_1157,net_1158})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'hAAAA"),
    .INIT_LUTF1("16'h0500"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_588
  (
    .clk(gclk_8),
    .ce(net_1165),
    .sr(net_182),
    .a({net_1302,net_1155}),
    .c({net_1182,open_n888}),
    .d({net_1312,open_n889}),
    .e({net_948,net_920}),
    .mi({open_n890,io_i2c_sda}),
    .f({net_1161,net_1165}),
    .q({open_n891,net_1166})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h5000"),
    .INIT_LUT1("16'h0400"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_589
  (
    .clk(gclk_8),
    .ce(net_1162),
    .sr(net_182),
    .a({net_1312,net_247}),
    .b({net_1182,open_n892}),
    .c({net_1302,net_1047}),
    .d({net_948,net_1155}),
    .mi({open_n893,io_i2c_sda}),
    .f({net_1155,net_1162}),
    .q({open_n894,net_1163})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0088"),
    .INIT_LUT1("16'h5505"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_590
  (
    .clk(gclk_8),
    .ce(net_1164),
    .sr(net_182),
    .a({net_960,net_961}),
    .b({open_n895,net_1047}),
    .c({net_961,open_n896}),
    .d({net_247,net_247}),
    .mi({open_n897,io_i2c_sda}),
    .f({net_1159,net_1164}),
    .q({open_n898,net_1167})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h000A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD_CARRY"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_591
  (
    .clk(gclk_9),
    .a({net_1461,1'b0}),
    .mi({open_n899,net_1461}),
    .f({net_1168,open_n900}),
    .q({open_n901,net_1173}),
    .fco(block_591_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_592
  (
    .clk(gclk_9),
    .a({net_1324,1'b0}),
    .b({1'b0,net_1460}),
    .mi({net_1324,net_1460}),
    .fci(block_591_carry),
    .f({net_1171,net_1169}),
    .q({net_1170,net_1172}),
    .fco(block_592_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_593
  (
    .clk(gclk_9),
    .a({1'b0,1'b0}),
    .b({net_1331,net_1198}),
    .mi({net_1331,net_1198}),
    .fci(block_592_carry),
    .f({net_1178,net_1179}),
    .q({net_1176,net_1175}),
    .fco(block_593_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_594
  (
    .clk(gclk_9),
    .a({net_1330,1'b0}),
    .b({1'b0,net_1203}),
    .mi({net_1330,net_1203}),
    .fci(block_593_carry),
    .f({net_1180,net_1174}),
    .q({net_1177,net_1181}),
    .fco(block_594_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_595
  (
    .clk(gclk_9),
    .a({1'b0,net_1202}),
    .b({net_1069,1'b0}),
    .mi({net_1069,net_1202}),
    .fci(block_594_carry),
    .f({net_1194,net_1185}),
    .q({net_1193,net_1187}),
    .fco(block_595_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_598
  (
    .clk(gclk_9),
    .a({net_1070,1'b0}),
    .b({1'b0,net_1075}),
    .mi({net_1075,net_1070}),
    .fci(block_595_carry),
    .f({net_1191,net_1188}),
    .q({net_1190,net_1195}),
    .fco(block_598_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_599
  (
    .clk(gclk_9),
    .a({open_n902,net_1074}),
    .b({open_n903,1'b0}),
    .mi({open_n904,net_1074}),
    .fci(block_598_carry),
    .f({open_n905,net_1196}),
    .q({open_n906,net_1197})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'hFEAA"),
    .INIT_LUTF1("16'hA888"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_596
  (
    .clk(gclk_8),
    .ce(net_1530),
    .sr(net_182),
    .a({net_967,net_1184}),
    .b({net_1300,net_1300}),
    .c({net_1532,net_1301}),
    .d({net_1301,net_1186}),
    .e({net_247,net_1299}),
    .mi({open_n907,net_1320}),
    .f({net_1184,net_1189}),
    .q({open_n908,net_1186})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hFFEE"),
    .INIT_LUTG0("16'hEF99"),
    .INIT_LUTF1("16'h00B0"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_597
  (
    .clk(gclk_8),
    .ce(net_1530),
    .sr(net_182),
    .a({net_1183,net_1182}),
    .b({net_1289,net_948}),
    .c({net_859,net_1078}),
    .d({net_1057,net_1302}),
    .e({net_1064,net_1312}),
    .mi({open_n909,net_1309}),
    .f({net_1192,net_1183}),
    .q({open_n910,net_1182})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0545"),
    .INIT_LUTG0("16'h5545"),
    .INIT_LUTF1("16'h0C0F"),
    .INIT_LUTG1("16'h0003"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("INV"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_600
  (
    .clk(gclk_9),
    .ce(i_mcu_dcs),
    .a({open_n911,net_1199}),
    .b({net_896,net_1198}),
    .c({i_mcu_rws,i_mcu_rws}),
    .d({net_1198,net_1142}),
    .e({net_1179,io_mcu_d[3]}),
    .f({net_1199,open_n912}),
    .q({open_n913,net_1198})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0503"),
    .INIT_LUT1("16'h0503"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_601
  (
    .a({net_1185,net_1196}),
    .b({net_1202,net_1074}),
    .c({i_mcu_rws,i_mcu_rws}),
    .d({net_896,net_896}),
    .f({net_1200,net_1201})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hCFAF"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("INV"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_602
  (
    .clk(gclk_9),
    .ce(i_mcu_dcs),
    .a({io_mcu_d[7],net_1202}),
    .b({net_1142,io_mcu_d[7]}),
    .c({i_mcu_rws,i_mcu_rws}),
    .d({net_1202,net_1142}),
    .mi({open_n914,net_1200}),
    .q({open_n915,net_1202})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0545"),
    .INIT_LUTG0("16'h5545"),
    .INIT_LUTF1("16'h000F"),
    .INIT_LUTG1("16'h0505"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("INV"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_603
  (
    .clk(gclk_9),
    .ce(i_mcu_dcs),
    .a({net_1174,net_1204}),
    .b({open_n916,net_1203}),
    .c({i_mcu_rws,i_mcu_rws}),
    .d({net_1203,net_1142}),
    .e({net_896,io_mcu_d[5]}),
    .f({net_1204,open_n917}),
    .q({open_n918,net_1203})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hBB0B"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_608
  (
    .a({net_974,net_1085}),
    .b({net_1085,net_974}),
    .c({net_1334,net_1334}),
    .d({net_1091,net_1091}),
    .mi({open_n919,net_1081}),
    .fx({open_n920,net_1208})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0045"),
    .INIT_LUTG0("16'h45FF"),
    .INIT_LUTF1("16'hF351"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_609
  (
    .a({net_881,net_1206}),
    .b({net_1085,net_1085}),
    .c({net_974,net_974}),
    .d({net_1205,net_1334}),
    .e({net_1082,net_1091}),
    .f({net_1206,net_1207})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hCCAA"),
    .INIT_LUT1("16'h0F0F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_610
  (
    .clk(gclk_4),
    .a({net_981,net_1205}),
    .b({net_994,net_981}),
    .c({net_511,net_511}),
    .d({net_1205,net_994}),
    .mi({open_n921,net_445}),
    .q({open_n922,net_1205})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hAFCF"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_611
  (
    .a({net_1545,net_1545}),
    .b({net_1538,net_1538}),
    .c({net_1044,net_189}),
    .d({net_189,net_1044}),
    .mi({open_n923,net_869}),
    .fx({open_n924,net_1209})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h00CF"),
    .INIT_LUTG0("16'h00AF"),
    .INIT_LUTF1("16'h1515"),
    .INIT_LUTG1("16'h0404"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_612
  (
    .clk(gclk_4),
    .a({net_189,net_1548}),
    .b({net_1044,net_1539}),
    .c({net_704,net_189}),
    .d({open_n925,net_1210}),
    .e({net_698,net_1044}),
    .mi({open_n926,net_1234}),
    .f({net_1210,net_1212}),
    .q({open_n927,net_1211})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h000A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD_CARRY"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("F"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_613
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1215,1'b0}),
    .q({net_1215,open_n928}),
    .fco(block_613_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_616
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1214,net_1216}),
    .b({1'b0,1'b0}),
    .fci(block_613_carry),
    .q({net_1214,net_1216}),
    .fco(block_616_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_617
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1224,net_1227}),
    .b({1'b0,1'b0}),
    .fci(block_616_carry),
    .q({net_1224,net_1227}),
    .fco(block_617_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_619
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1223,net_1226}),
    .b({1'b0,1'b0}),
    .fci(block_617_carry),
    .q({net_1223,net_1226}),
    .fco(block_619_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_620
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1232,net_1234}),
    .b({1'b0,1'b0}),
    .fci(block_619_carry),
    .q({net_1232,net_1234}),
    .fco(block_620_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_621
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1231,net_1233}),
    .b({1'b0,1'b0}),
    .fci(block_620_carry),
    .q({net_1231,net_1233}),
    .fco(block_621_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_623
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({open_n929,net_1241}),
    .b({open_n930,1'b0}),
    .fci(block_621_carry),
    .q({open_n931,net_1241})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h7771"),
    .INIT_LUTF1("16'hA800"),
    .INIT_LUTG1("16'hAAA8"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_614
  (
    .clk(gclk_9),
    .ce(net_882),
    .a({net_1343,net_1213}),
    .b({net_1090,net_623}),
    .c({net_1098,net_1088}),
    .d({net_1213,net_1089}),
    .e({net_623,net_1344}),
    .mi({open_n932,io_mcu_d[7]}),
    .f({net_1221,net_1220}),
    .q({open_n933,net_1213})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'hAAA8"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hFBFB"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_615
  (
    .clk(gclk_4),
    .a({net_1215,net_1231}),
    .b({net_1105,net_1234}),
    .c({net_1216,net_1232}),
    .d({open_n934,net_1217}),
    .e({net_1223,net_1233}),
    .mi({net_1215,net_1231}),
    .f({net_1217,net_1222}),
    .q({net_1219,net_1218})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hF3B2"),
    .INIT_LUTG0("16'hB230"),
    .INIT_LUTF1("16'hFF55"),
    .INIT_LUTG1("16'hF550"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_618
  (
    .clk(gclk_9),
    .ce(net_897),
    .a({net_1225,net_1228}),
    .b({open_n935,net_899}),
    .c({net_1352,net_1359}),
    .d({net_1353,net_1351}),
    .e({net_898,net_1230}),
    .mi({io_mcu_d[1],io_mcu_d[2]}),
    .f({net_1228,net_1229}),
    .q({net_1225,net_1230})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h7700"),
    .INIT_LUTG0("16'h0700"),
    .INIT_LUTF1("16'h3F3F"),
    .INIT_LUTG1("16'h1515"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_622
  (
    .clk(gclk_4),
    .a({net_1251,net_906}),
    .b({i_adc2B_d[5],net_1043}),
    .c({net_1242,i_adc1A_d[5]}),
    .d({open_n936,net_1235}),
    .e({i_adc2A_d[5],net_1244}),
    .mi({i_adc2A_d[5],i_adc1A_d[5]}),
    .f({net_1235,net_1238}),
    .q({net_1236,net_1237})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h135F"),
    .INIT_LUTF1("16'h0700"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_624
  (
    .clk(gclk_4),
    .a({net_1244,net_1242}),
    .b({i_adc1A_d[2],i_adc2A_d[2]}),
    .c({net_1125,i_adc2B_d[2]}),
    .d({net_1240,net_1251}),
    .e({net_1513,net_1017}),
    .mi({i_adc1A_d[2],i_adc2A_d[2]}),
    .f({net_1247,net_1240}),
    .q({net_1250,net_1248})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h1000"),
    .INIT_LUT1("16'h8000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_625
  (
    .clk(gclk_4),
    .a({net_308,net_180}),
    .b({net_181,net_181}),
    .c({net_180,net_308}),
    .d({net_536,net_536}),
    .mi({i_adc2B_d[5],i_adc2B_d[0]}),
    .f({net_1242,net_1244}),
    .q({net_1243,net_1246})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0101"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hF0F0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_626
  (
    .clk(gclk_0),
    .sr(net_1498),
    .a({open_n937,net_1239}),
    .b({open_n938,net_1356}),
    .c({net_1500,net_1255}),
    .e({net_823,net_1360}),
    .mi({open_n939,net_1366}),
    .f({net_1245,net_1249}),
    .q({open_n940,net_1239})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0777"),
    .INIT_LUT1("16'h8888"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_627
  (
    .clk(gclk_4),
    .a({net_249,net_794}),
    .b({net_536,i_adc1B_d[0]}),
    .c({open_n941,i_adc2A_d[0]}),
    .d({open_n942,net_1251}),
    .mi({i_adc2B_d[2],i_adc2A_d[0]}),
    .f({net_1251,net_1258}),
    .q({net_1254,net_1257})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0002"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0001"),
    .INIT_LUTG1("16'h0001"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_628
  (
    .clk(gclk_0),
    .sr(net_1498),
    .a({net_1357,net_1252}),
    .b({net_1363,net_1497}),
    .c({net_1381,net_1256}),
    .d({net_1369,net_1382}),
    .e({open_n943,net_1372}),
    .mi({net_1365,net_1374}),
    .f({net_1252,net_1253}),
    .q({net_1255,net_1256})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hAAFF"),
    .INIT_LUTG0("16'h303F"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h1000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_629
  (
    .clk(gclk_9),
    .ce(net_1259),
    .a({net_1264,net_778}),
    .b({net_1508,net_1264}),
    .c({net_1263,net_632}),
    .d({net_1145,net_1127}),
    .e({net_1507,i_mcu_rws}),
    .mi({io_mcu_d[0],io_mcu_d[5]}),
    .f({net_1259,net_1262}),
    .q({net_1260,net_1261})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h000A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD_CARRY"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("F"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_630
  (
    .clk(gclk_4),
    .ce(net_994),
    .sr(net_445),
    .a({net_1266,1'b0}),
    .q({net_1266,open_n944}),
    .fco(block_630_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_633
  (
    .clk(gclk_4),
    .ce(net_994),
    .sr(net_445),
    .a({net_1265,net_1267}),
    .b({1'b0,1'b0}),
    .fci(block_630_carry),
    .q({net_1265,net_1267}),
    .fco(block_633_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_634
  (
    .clk(gclk_4),
    .ce(net_994),
    .sr(net_445),
    .a({net_1273,net_1275}),
    .b({1'b0,1'b0}),
    .fci(block_633_carry),
    .q({net_1273,net_1275}),
    .fco(block_634_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_636
  (
    .clk(gclk_4),
    .ce(net_994),
    .sr(net_445),
    .a({net_1272,net_1274}),
    .b({1'b0,1'b0}),
    .fci(block_634_carry),
    .q({net_1272,net_1274}),
    .fco(block_636_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_637
  (
    .clk(gclk_4),
    .ce(net_994),
    .sr(net_445),
    .a({net_1280,net_1282}),
    .b({1'b0,1'b0}),
    .fci(block_636_carry),
    .q({net_1280,net_1282}),
    .fco(block_637_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_638
  (
    .clk(gclk_4),
    .ce(net_994),
    .sr(net_445),
    .a({net_1279,net_1281}),
    .b({1'b0,1'b0}),
    .fci(block_637_carry),
    .q({net_1279,net_1281}),
    .fco(block_638_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_640
  (
    .clk(gclk_4),
    .ce(net_994),
    .sr(net_445),
    .a({open_n945,net_1288}),
    .b({open_n946,1'b0}),
    .fci(block_638_carry),
    .q({open_n947,net_1288})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0A33"),
    .INIT_LUTG0("16'h0A3B"),
    .INIT_LUTF1("16'h0A33"),
    .INIT_LUTG1("16'h0A3B"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_631
  (
    .clk(gclk_9),
    .a({net_1263,net_1264}),
    .b({net_1268,net_1262}),
    .c({i_mcu_rws,i_mcu_rws}),
    .d({i_mcu_dcs,i_mcu_dcs}),
    .e({net_778,net_778}),
    .q({net_1263,net_1264})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hAAFF"),
    .INIT_LUTG0("16'h303F"),
    .INIT_LUTF1("16'h0400"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_632
  (
    .clk(gclk_9),
    .ce(net_1269),
    .a({net_1507,net_778}),
    .b({net_1263,net_1263}),
    .c({net_1264,net_632}),
    .d({net_1145,net_1128}),
    .e({net_1508,i_mcu_rws}),
    .mi({io_mcu_d[2],io_mcu_d[1]}),
    .f({net_1269,net_1268}),
    .q({net_1270,net_1271})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h2222"),
    .INIT_LUTF1("16'h0004"),
    .INIT_LUTG1("16'h0004"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_635
  (
    .clk(gclk_8),
    .ce(net_1277),
    .sr(net_182),
    .a({net_1301,net_1276}),
    .b({net_1300,net_247}),
    .c({net_1299,open_n948}),
    .d({net_1532,open_n949}),
    .e({open_n950,net_1521}),
    .mi({open_n951,io_i2c_sda}),
    .f({net_1276,net_1277}),
    .q({open_n952,net_1278})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0003"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0044"),
    .INIT_LUTG1("16'h00CC"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_639
  (
    .clk(gclk_9),
    .ce(net_1156),
    .a({net_1283,open_n953}),
    .b({net_439,net_1263}),
    .c({open_n954,net_1507}),
    .d({net_1034,net_1508}),
    .e({net_1292,net_1264}),
    .mi({io_mcu_d[2],io_mcu_d[1]}),
    .f({net_1286,net_1283}),
    .q({net_1284,net_1285})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hFC30"),
    .INIT_LUTG0("16'hFC30"),
    .INIT_LUTF1("16'h0F0F"),
    .INIT_LUTG1("16'h0F0F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_641
  (
    .clk(gclk_4),
    .ce(net_1291),
    .sr(net_445),
    .b({open_n955,net_527}),
    .c({net_1348,net_1281}),
    .d({open_n956,net_1190}),
    .mi({net_1266,net_1281}),
    .f({net_1291,net_1294}),
    .q({net_1297,net_1296})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0001"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h0001"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_642
  (
    .clk(gclk_8),
    .ce(net_1530),
    .sr(net_182),
    .a({net_1314,net_1287}),
    .b({net_1311,net_1311}),
    .c({net_1186,net_1314}),
    .d({net_1287,net_1062}),
    .e({net_1531,net_1531}),
    .mi({open_n957,net_1316}),
    .f({net_1289,net_1295}),
    .q({open_n958,net_1287})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hFA0A"),
    .INIT_LUT1("16'hFC0C"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_643
  (
    .clk(gclk_4),
    .ce(net_1291),
    .sr(net_445),
    .a({open_n959,net_1280}),
    .b({net_1267,open_n960}),
    .c({net_527,net_527}),
    .d({net_1172,net_1193}),
    .mi({net_1267,net_1280}),
    .f({net_1290,net_1298}),
    .q({net_1293,net_1292})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h000A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_644
  (
    .clk(gclk_8),
    .ce(net_1530),
    .sr(net_182),
    .a({net_1301,1'b0}),
    .b({net_1300,net_1532}),
    .c({1'b0,1'b0}),
    .d({1'b0,open_n961}),
    .e({1'b0,open_n962}),
    .mi({net_1304,net_1305}),
    .f({net_1305,open_n963}),
    .fx({net_1304,net_1308}),
    .q({net_1300,net_1301}),
    .fco(sig_644_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_645
  (
    .clk(gclk_8),
    .ce(net_1530),
    .sr(net_182),
    .a({net_948,net_1299}),
    .b({net_1182,net_1302}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1306,net_1307}),
    .fci(sig_644_carry),
    .f({net_1310,net_1307}),
    .fx({net_1309,net_1306}),
    .q({net_1302,net_1299}),
    .fco(sig_645_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_647
  (
    .clk(gclk_8),
    .ce(net_1530),
    .sr(net_182),
    .a({net_1287,net_1312}),
    .b({net_1314,net_1186}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1318,net_1322}),
    .fci(sig_645_carry),
    .f({net_1316,net_1318}),
    .fx({net_1322,net_1320}),
    .q({net_1312,net_1314}),
    .fco(sig_647_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_648
  (
    .clk(gclk_8),
    .ce(net_1530),
    .sr(net_182),
    .a({net_1325,net_1311}),
    .b({net_1529,net_1313}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1317,net_1321}),
    .fci(sig_647_carry),
    .f({net_1319,net_1321}),
    .fx({net_1315,net_1317}),
    .q({net_1313,net_1311}),
    .fco(sig_648_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_649
  (
    .clk(gclk_8),
    .ce(net_1530),
    .sr(net_182),
    .a({open_n964,net_1323}),
    .c({1'b0,1'b0}),
    .d({open_n965,1'b0}),
    .mi({open_n966,net_1328}),
    .fci(sig_648_carry),
    .f({open_n967,net_1328}),
    .q({open_n968,net_1323})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h0400"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_646
  (
    .a({net_1301,net_1301}),
    .b({net_1289,net_1532}),
    .c({net_1532,net_1289}),
    .d({net_1300,net_1300}),
    .mi({open_n969,net_1299}),
    .fx({open_n970,net_1303})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h00AF"),
    .INIT_LUTG0("16'h00CF"),
    .INIT_LUTF1("16'h0033"),
    .INIT_LUTG1("16'h0303"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("INV"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_650
  (
    .clk(gclk_9),
    .ce(i_mcu_dcs),
    .a({open_n971,net_1324}),
    .b({i_mcu_rws,io_mcu_d[2]}),
    .c({net_1171,i_mcu_rws}),
    .d({net_1324,net_1326}),
    .e({net_896,net_1142}),
    .f({net_1326,open_n972}),
    .q({open_n973,net_1324})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hAAA8"),
    .INIT_LUT1("16'h1000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_651
  (
    .clk(gclk_8),
    .ce(net_1530),
    .sr(net_182),
    .a({net_1182,net_1325}),
    .b({net_948,net_1052}),
    .c({net_1312,net_1311}),
    .d({net_1302,net_1313}),
    .mi({open_n974,net_1319}),
    .f({net_1329,net_1327}),
    .q({open_n975,net_1325})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hCFAF"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("INV"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_652
  (
    .clk(gclk_9),
    .ce(i_mcu_dcs),
    .a({io_mcu_d[6],net_1330}),
    .b({net_1142,io_mcu_d[6]}),
    .c({i_mcu_rws,i_mcu_rws}),
    .d({net_1330,net_1142}),
    .mi({open_n976,net_1033}),
    .q({open_n977,net_1330})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0545"),
    .INIT_LUTG0("16'h5545"),
    .INIT_LUTF1("16'h0033"),
    .INIT_LUTG1("16'h1111"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("INV"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_653
  (
    .clk(gclk_9),
    .ce(i_mcu_dcs),
    .a({net_1178,net_1332}),
    .b({i_mcu_rws,net_1331}),
    .c({open_n978,i_mcu_rws}),
    .d({net_1331,net_1142}),
    .e({net_896,io_mcu_d[4]}),
    .f({net_1332,open_n979}),
    .q({open_n980,net_1331})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h2000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_654
  (
    .a({net_1182,net_1312}),
    .b({net_1312,net_1302}),
    .c({net_948,net_948}),
    .d({net_1302,net_1182}),
    .mi({open_n981,net_1289}),
    .fx({open_n982,net_1333})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hCCAA"),
    .INIT_LUT1("16'h0F0F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_655
  (
    .clk(gclk_4),
    .a({net_1084,net_1334}),
    .b({net_994,net_1084}),
    .c({net_511,net_511}),
    .d({net_1334,net_994}),
    .mi({open_n983,net_445}),
    .q({open_n984,net_1334})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA220"),
    .INIT_LUTG0("16'hA2A2"),
    .INIT_LUTF1("16'h50D0"),
    .INIT_LUTG1("16'hD0F0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_656
  (
    .a({net_1094,net_1094}),
    .b({net_1207,net_1079}),
    .c({net_1342,net_1086}),
    .d({net_1079,net_1477}),
    .e({net_1086,net_1208}),
    .f({net_1336,net_1335})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h5555"),
    .INIT_LUT1("16'hFFCF"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_657
  (
    .clk(gclk_2),
    .ce(net_1338),
    .a({open_n985,net_1337}),
    .b({net_1481,open_n986}),
    .c({net_1476,open_n987}),
    .d({net_1473,open_n988}),
    .f({net_1338,open_n989}),
    .q({open_n990,net_1337})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h4455"),
    .INIT_LUTG0("16'h4054"),
    .INIT_LUTF1("16'h0045"),
    .INIT_LUTG1("16'h4555"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_658
  (
    .a({net_1350,net_1350}),
    .b({net_1092,net_875}),
    .c({net_1482,net_1482}),
    .d({net_875,net_1213}),
    .e({net_1213,net_1092}),
    .f({net_1342,net_1339})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0100"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h0777"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_659
  (
    .clk(gclk_4),
    .a({net_1251,net_794}),
    .b({i_adc2A_d[3],net_1251}),
    .c({net_1242,net_1242}),
    .d({i_adc2B_d[3],net_649}),
    .e({net_1021,net_778}),
    .mi({i_adc2A_d[3],i_adc2B_d[3]}),
    .f({net_1345,net_1341}),
    .q({net_1340,net_1346})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h3311"),
    .INIT_LUT1("16'h2222"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_660
  (
    .a({net_511,net_1339}),
    .b({net_1336,net_511}),
    .d({open_n991,net_1335}),
    .f({net_1343,net_1344})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h5555"),
    .INIT_LUTG0("16'h5555"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'hF0F0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_661
  (
    .clk(gclk_5),
    .ce(net_1665),
    .a({open_n992,net_1347}),
    .c({net_309,open_n993}),
    .e({net_249,open_n994}),
    .f({net_1349,open_n995}),
    .q({open_n996,net_1347})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hFFEE"),
    .INIT_LUTG0("16'hFFEE"),
    .INIT_LUTF1("16'hF0F0"),
    .INIT_LUTG1("16'hFFFF"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_662
  (
    .clk(gclk_4),
    .ce(net_1140),
    .sr(net_445),
    .a({open_n997,net_1348}),
    .b({open_n998,net_1220}),
    .c({net_1344,open_n999}),
    .d({open_n1000,net_1221}),
    .e({net_1343,open_n1001}),
    .q({net_1350,net_1348})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h000A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD_CARRY"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("F"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_663
  (
    .clk(gclk_6),
    .sr(net_1112),
    .a({net_1352,1'b0}),
    .q({net_1352,open_n1002}),
    .fco(block_663_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_664
  (
    .clk(gclk_6),
    .sr(net_1112),
    .a({net_1351,net_1353}),
    .b({1'b0,1'b0}),
    .fci(block_663_carry),
    .q({net_1351,net_1353}),
    .fco(block_664_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_665
  (
    .clk(gclk_6),
    .sr(net_1112),
    .a({net_1355,net_1359}),
    .b({1'b0,1'b0}),
    .fci(block_664_carry),
    .q({net_1355,net_1359}),
    .fco(block_665_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_667
  (
    .clk(gclk_6),
    .sr(net_1112),
    .a({net_1354,net_1358}),
    .b({1'b0,1'b0}),
    .fci(block_665_carry),
    .q({net_1354,net_1358}),
    .fco(block_667_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_669
  (
    .clk(gclk_6),
    .sr(net_1112),
    .a({open_n1003,net_1370}),
    .b({open_n1004,1'b0}),
    .fci(block_667_carry),
    .q({open_n1005,net_1370})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h000A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_666
  (
    .clk(gclk_0),
    .sr(net_1498),
    .a({net_1357,1'b0}),
    .b({net_1239,net_1363}),
    .c({1'b0,1'b0}),
    .d({1'b0,open_n1006}),
    .e({1'b0,open_n1007}),
    .mi({net_1361,net_1368}),
    .f({net_1361,open_n1008}),
    .fx({net_1366,net_1368}),
    .q({net_1357,net_1363}),
    .fco(sig_666_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_668
  (
    .clk(gclk_0),
    .sr(net_1498),
    .a({net_1255,net_1356}),
    .b({net_1493,net_1360}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1364,net_1367}),
    .fci(sig_666_carry),
    .f({net_1365,net_1367}),
    .fx({net_1362,net_1364}),
    .q({net_1360,net_1356}),
    .fco(sig_668_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_670
  (
    .clk(gclk_0),
    .sr(net_1498),
    .a({net_1494,net_1371}),
    .b({net_1381,net_1385}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1376,net_1380}),
    .fci(sig_668_carry),
    .f({net_1373,net_1376}),
    .fx({net_1380,net_1378}),
    .q({net_1371,net_1381}),
    .fco(sig_670_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_671
  (
    .clk(gclk_0),
    .sr(net_1498),
    .a({net_1497,net_1369}),
    .b({net_1256,net_1372}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1375,net_1379}),
    .fci(sig_670_carry),
    .f({net_1377,net_1379}),
    .fx({net_1374,net_1375}),
    .q({net_1372,net_1369}),
    .fco(sig_671_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_673
  (
    .clk(gclk_0),
    .sr(net_1498),
    .a({open_n1009,net_1382}),
    .c({1'b0,1'b0}),
    .d({open_n1010,1'b0}),
    .mi({net_1378,net_1384}),
    .fci(sig_671_carry),
    .f({open_n1011,net_1384}),
    .q({net_1385,net_1382})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h000A"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB_CARRY"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_672
  (
    .a({net_1260,1'b0}),
    .b({net_1396,open_n1012}),
    .fco(block_672_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_674
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1124,net_1123}),
    .b({net_1383,net_1395}),
    .mi({open_n1013,net_1398}),
    .fci(block_672_carry),
    .q({open_n1014,net_1383}),
    .fco(block_674_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_675
  (
    .clk(gclk_9),
    .ce(net_1259),
    .a({net_1386,net_1387}),
    .b({net_1397,net_1394}),
    .mi({io_mcu_d[4],io_mcu_d[3]}),
    .fci(block_674_carry),
    .q({net_1386,net_1387}),
    .fco(block_675_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_677
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1138,net_1261}),
    .b({net_1388,net_1391}),
    .mi({net_1401,net_1404}),
    .fci(block_675_carry),
    .q({net_1388,net_1391}),
    .fco(block_677_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_678
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1393,net_1137}),
    .b({net_1403,net_1413}),
    .mi({open_n1015,net_1415}),
    .fci(block_677_carry),
    .q({open_n1016,net_1403}),
    .fco(block_678_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_681
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1270,net_1271}),
    .b({net_1412,net_1400}),
    .mi({open_n1017,net_1414}),
    .fci(block_678_carry),
    .q({open_n1018,net_1400}),
    .fco(block_681_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_682
  (
    .clk(gclk_9),
    .ce(net_1269),
    .a({net_1407,net_1409}),
    .b({net_1422,net_1408}),
    .mi({io_mcu_d[4],io_mcu_d[3]}),
    .fci(block_681_carry),
    .q({net_1407,net_1409}),
    .fco(block_682_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_685
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1143,net_1389}),
    .b({net_1410,net_1411}),
    .mi({net_1416,net_1419}),
    .fci(block_682_carry),
    .q({net_1410,net_1411}),
    .fco(block_685_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_686
  (
    .clk(gclk_9),
    .ce(net_1269),
    .a({net_1151,net_1425}),
    .b({net_1434,net_1423}),
    .mi({open_n1019,io_mcu_d[7]}),
    .fci(block_685_carry),
    .q({open_n1020,net_1425}),
    .fco(block_686_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_689
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1039,net_1153}),
    .b({net_1432,net_1429}),
    .mi({net_1428,net_1433}),
    .fci(block_686_carry),
    .q({net_1432,net_1429}),
    .fco(block_689_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_690
  (
    .clk(gclk_9),
    .ce(net_1149),
    .a({net_1439,net_1441}),
    .b({net_1427,net_1424}),
    .mi({io_mcu_d[4],io_mcu_d[3]}),
    .fci(block_689_carry),
    .q({net_1439,net_1441}),
    .fco(block_690_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_693
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_917,net_1037}),
    .b({net_1449,net_1446}),
    .mi({net_1431,net_1426}),
    .fci(block_690_carry),
    .q({net_1449,net_1446}),
    .fco(block_693_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_694
  (
    .clk(gclk_9),
    .ce(net_1149),
    .a({net_1157,net_1455}),
    .b({net_1443,net_1438}),
    .mi({open_n1021,io_mcu_d[7]}),
    .fci(block_693_carry),
    .q({open_n1022,net_1455}),
    .fco(block_694_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_696
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1284,net_1285}),
    .b({net_1456,net_1458}),
    .mi({net_1445,net_1447}),
    .fci(block_694_carry),
    .q({net_1456,net_1458}),
    .fco(block_696_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_697
  (
    .clk(gclk_9),
    .ce(net_1156),
    .a({net_1459,net_1462}),
    .b({net_1444,net_1440}),
    .mi({io_mcu_d[4],io_mcu_d[3]}),
    .fci(block_696_carry),
    .q({net_1459,net_1462}),
    .fco(block_697_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_700
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1019,net_1158}),
    .b({net_1465,net_1466}),
    .mi({net_1450,net_1442}),
    .fci(block_697_carry),
    .q({net_1465,net_1466}),
    .fco(block_700_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h999C"),
    .INIT_LUT1("16'h999C"),
    .ALUTYPE("SUB"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_701
  (
    .clk(gclk_9),
    .ce(net_1156),
    .a({1'b0,net_1467}),
    .b({open_n1023,net_1454}),
    .mi({open_n1024,io_mcu_d[7]}),
    .fci(block_700_carry),
    .f({net_1469,open_n1025}),
    .q({open_n1026,net_1467})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hAAFF"),
    .INIT_LUTG0("16'h303F"),
    .INIT_LUTF1("16'hAFAF"),
    .INIT_LUTG1("16'h330F"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_676
  (
    .clk(gclk_9),
    .ce(net_1269),
    .a({net_778,net_778}),
    .b({net_1507,net_1508}),
    .c({net_1129,net_632}),
    .d({net_632,net_1132}),
    .e({i_mcu_rws,i_mcu_rws}),
    .mi({io_mcu_d[5],io_mcu_d[0]}),
    .f({net_1390,net_1392}),
    .q({net_1389,net_1393})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h000A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_679
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1395,1'b0}),
    .b({net_1383,net_1396}),
    .c({1'b0,1'b0}),
    .d({1'b0,open_n1027}),
    .e({1'b0,open_n1028}),
    .mi({net_1399,net_1405}),
    .f({net_1399,open_n1029}),
    .fx({net_1398,net_1405}),
    .q({net_1395,net_1396}),
    .fco(sig_679_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_680
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1391,net_1394}),
    .b({net_1388,net_1397}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1402,net_1406}),
    .fci(sig_679_carry),
    .f({net_1404,net_1406}),
    .fx({net_1401,net_1402}),
    .q({net_1397,net_1394}),
    .fco(sig_680_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_683
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1400,net_1413}),
    .b({net_1412,net_1403}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1418,net_1421}),
    .fci(sig_680_carry),
    .f({net_1414,net_1418}),
    .fx({net_1421,net_1415}),
    .q({net_1413,net_1412}),
    .fco(sig_683_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_684
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1411,net_1408}),
    .b({net_1410,net_1422}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1417,net_1420}),
    .fci(sig_683_carry),
    .f({net_1419,net_1420}),
    .fx({net_1416,net_1417}),
    .q({net_1422,net_1408}),
    .fco(sig_684_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_687
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1429,net_1423}),
    .b({net_1432,net_1434}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1436,net_1430}),
    .fci(sig_684_carry),
    .f({net_1433,net_1430}),
    .fx({net_1428,net_1436}),
    .q({net_1434,net_1423}),
    .fco(sig_687_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_688
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1446,net_1424}),
    .b({net_1449,net_1427}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1435,net_1437}),
    .fci(sig_687_carry),
    .f({net_1426,net_1437}),
    .fx({net_1431,net_1435}),
    .q({net_1427,net_1424}),
    .fco(sig_688_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_691
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1458,net_1438}),
    .b({net_1456,net_1443}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1452,net_1448}),
    .fci(sig_688_carry),
    .f({net_1447,net_1448}),
    .fx({net_1445,net_1452}),
    .q({net_1443,net_1438}),
    .fco(sig_691_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_692
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({net_1466,net_1440}),
    .b({net_1465,net_1444}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1451,net_1453}),
    .fci(sig_691_carry),
    .f({net_1442,net_1453}),
    .fx({net_1450,net_1451}),
    .q({net_1444,net_1440}),
    .fco(sig_692_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_695
  (
    .clk(gclk_4),
    .sr(net_445),
    .a({open_n1030,net_1454}),
    .c({1'b0,1'b0}),
    .d({open_n1031,1'b0}),
    .mi({open_n1032,net_1457}),
    .fci(sig_692_carry),
    .f({open_n1033,net_1457}),
    .q({open_n1034,net_1454})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0545"),
    .INIT_LUTG0("16'h5545"),
    .INIT_LUTF1("16'h4477"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("INV"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_698
  (
    .clk(gclk_9),
    .ce(i_mcu_dcs),
    .a({net_1168,net_1464}),
    .b({net_896,net_1461}),
    .c({open_n1035,i_mcu_rws}),
    .d({net_1461,net_1142}),
    .e({i_mcu_rws,io_mcu_d[0]}),
    .f({net_1464,open_n1036}),
    .q({open_n1037,net_1461})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h00AF"),
    .INIT_LUTG0("16'h00CF"),
    .INIT_LUTF1("16'h4477"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("INV"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_699
  (
    .clk(gclk_9),
    .ce(i_mcu_dcs),
    .a({net_1169,net_1460}),
    .b({net_896,io_mcu_d[1]}),
    .c({open_n1038,i_mcu_rws}),
    .d({net_1460,net_1463}),
    .e({i_mcu_rws,net_1142}),
    .f({net_1463,open_n1039}),
    .q({open_n1040,net_1460})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h0020"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_702
  (
    .a({net_1182,net_948}),
    .b({net_948,net_1312}),
    .c({net_1289,net_1289}),
    .d({net_1312,net_1182}),
    .mi({open_n1041,net_1302}),
    .fx({open_n1042,net_1468})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hFFFF"),
    .INIT_LUTG0("16'hFF00"),
    .INIT_LUTF1("16'h5555"),
    .INIT_LUTG1("16'h5555"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_707
  (
    .clk(gclk_0),
    .ce(net_451),
    .a({net_1471,open_n1043}),
    .d({open_n1044,net_1471}),
    .e({open_n1045,net_901}),
    .q({net_1471,net_1472})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h000A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD_CARRY"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("F"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_708
  (
    .clk(gclk_2),
    .sr(net_1338),
    .a({net_1474,1'b0}),
    .q({net_1474,open_n1046}),
    .fco(block_708_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_710
  (
    .clk(gclk_2),
    .sr(net_1338),
    .a({net_1473,net_1475}),
    .b({1'b0,1'b0}),
    .fci(block_708_carry),
    .q({net_1473,net_1475}),
    .fco(block_710_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_711
  (
    .clk(gclk_2),
    .sr(net_1338),
    .a({net_1479,net_1481}),
    .b({1'b0,1'b0}),
    .fci(block_710_carry),
    .q({net_1479,net_1481}),
    .fco(block_711_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_712
  (
    .clk(gclk_2),
    .sr(net_1338),
    .a({net_1478,net_1480}),
    .b({1'b0,1'b0}),
    .fci(block_711_carry),
    .q({net_1478,net_1480}),
    .fco(block_712_carry)
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h666A"),
    .INIT_LUT1("16'h666A"),
    .ALUTYPE("ADD"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_713
  (
    .clk(gclk_2),
    .sr(net_1338),
    .a({open_n1047,net_1483}),
    .b({open_n1048,1'b0}),
    .fci(block_712_carry),
    .q({open_n1049,net_1483})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0003"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h5050"),
    .INIT_LUTG1("16'h5050"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_709
  (
    .a({net_1334,open_n1050}),
    .b({open_n1051,net_1480}),
    .c({net_1091,net_1478}),
    .d({open_n1052,net_1483}),
    .e({open_n1053,net_1479}),
    .f({net_1477,net_1476})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0AAA"),
    .INIT_LUTG0("16'h0222"),
    .INIT_LUTF1("16'h7777"),
    .INIT_LUTG1("16'h0707"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_714
  (
    .clk(gclk_4),
    .a({net_998,net_1485}),
    .b({net_827,i_adc2A_d[7]}),
    .c({net_999,i_adc2B_d[7]}),
    .d({open_n1054,net_1242}),
    .e({net_1278,net_1251}),
    .mi({i_adc2B_d[7],i_adc2A_d[7]}),
    .f({net_1485,net_1490}),
    .q({net_1488,net_1489})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h7700"),
    .INIT_LUTG0("16'h0700"),
    .INIT_LUTF1("16'h7777"),
    .INIT_LUTG1("16'h0707"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_715
  (
    .clk(gclk_4),
    .a({net_1042,net_1251}),
    .b({net_998,i_adc2A_d[4]}),
    .c({net_1242,net_999}),
    .d({open_n1055,net_1484}),
    .e({i_adc2B_d[4],net_1163}),
    .mi({i_adc2B_d[4],i_adc2A_d[4]}),
    .f({net_1484,net_1491}),
    .q({net_1486,net_1487})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hCCAA"),
    .INIT_LUT1("16'h3333"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("FX"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_716
  (
    .clk(gclk_4),
    .a({net_1100,net_1482}),
    .b({net_511,net_1100}),
    .c({net_994,net_511}),
    .d({net_1482,net_994}),
    .mi({open_n1056,net_445}),
    .q({open_n1057,net_1482})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h5555"),
    .INIT_LUTG0("16'h5555"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_717
  (
    .clk(gclk_0),
    .ce(net_1498),
    .a({open_n1058,net_1492}),
    .q({open_n1059,net_1492})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h2233"),
    .INIT_LUT1("16'hFC0C"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("INV"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_718
  (
    .clk(gclk_4),
    .ce(net_1499),
    .sr(net_445),
    .a({open_n1060,net_1115}),
    .b({net_1617,net_1348}),
    .c({net_527,open_n1061}),
    .d({i_mcu_clk,net_1469}),
    .mi({open_n1062,1'b0}),
    .f({net_1501,net_1499}),
    .q({open_n1063,net_1496})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0001"),
    .INIT_LUTF1("16'h33FF"),
    .INIT_LUTG1("16'h33FF"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_719
  (
    .clk(gclk_0),
    .sr(net_1498),
    .a({open_n1064,net_1493}),
    .b({net_1253,net_1494}),
    .c({open_n1065,net_1385}),
    .d({net_1495,net_1371}),
    .e({open_n1066,net_1249}),
    .mi({net_1377,net_1362}),
    .f({net_1498,net_1495}),
    .q({net_1497,net_1493})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'hBBBB"),
    .INIT_LUT1("16'h8800"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_720
  (
    .clk(gclk_0),
    .ce(net_451),
    .a({net_1648,net_1618}),
    .b({net_1289,net_901}),
    .d({net_952,open_n1067}),
    .f({net_1500,open_n1068}),
    .q({open_n1069,net_1502})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_721
  (
    .clk(gclk_0),
    .sr(net_1498),
    .mi({open_n1070,net_1373}),
    .q({open_n1071,net_1494})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h020A"),
    .INIT_LUTF1("16'h55FF"),
    .INIT_LUTG1("16'h1133"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_722
  (
    .clk(gclk_4),
    .a({net_998,net_1503}),
    .b({net_1251,i_adc2B_d[6]}),
    .c({open_n1072,net_1148}),
    .d({net_1522,net_1242}),
    .e({i_adc2A_d[6],net_1026}),
    .mi({i_adc2A_d[6],i_adc2B_d[6]}),
    .f({net_1503,net_1505}),
    .q({net_1504,net_1506})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0A33"),
    .INIT_LUTG0("16'h0A3B"),
    .INIT_LUTF1("16'h0AFF"),
    .INIT_LUTG1("16'h0A08"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_723
  (
    .clk(gclk_9),
    .a({net_1507,net_1508}),
    .b({net_778,net_1392}),
    .c({i_mcu_rws,i_mcu_rws}),
    .d({i_mcu_dcs,i_mcu_dcs}),
    .e({net_1390,net_778}),
    .q({net_1507,net_1508})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0808"),
    .INIT_LUT1("16'h30F0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_724
  (
    .clk(gclk_8),
    .ce(net_1514),
    .sr(net_182),
    .a({open_n1073,net_1276}),
    .b({net_796,net_584}),
    .c({net_1135,net_247}),
    .d({net_1509,open_n1074}),
    .mi({open_n1075,io_i2c_sda}),
    .f({net_1515,net_1514}),
    .q({open_n1076,net_1509})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hACAC"),
    .INIT_LUTG0("16'hACAC"),
    .INIT_LUTF1("16'hF000"),
    .INIT_LUTG1("16'hF000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("0"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_725
  (
    .clk(gclk_4),
    .a({open_n1077,net_1173}),
    .b({open_n1078,net_1266}),
    .c({i_adc1B_d[2],net_527}),
    .d({net_794,open_n1079}),
    .mi({i_adc1B_d[2],net_1216}),
    .f({net_1513,net_1512}),
    .q({net_1517,net_1511})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h00CC"),
    .INIT_LUTF1("16'h7777"),
    .INIT_LUTG1("16'h0077"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_726
  (
    .clk(gclk_8),
    .ce(net_1516),
    .sr(net_182),
    .a({net_999,open_n1080}),
    .b({net_1059,net_1276}),
    .d({net_1510,net_247}),
    .e({net_998,net_1523}),
    .mi({open_n1081,io_i2c_sda}),
    .f({net_1518,net_1516}),
    .q({open_n1082,net_1510})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0088"),
    .INIT_LUT1("16'hA0A0"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_727
  (
    .clk(gclk_8),
    .ce(net_1520),
    .sr(net_182),
    .a({net_1155,net_1155}),
    .b({open_n1083,net_1303}),
    .c({net_1289,open_n1084}),
    .d({open_n1085,net_247}),
    .mi({open_n1086,io_i2c_sda}),
    .f({net_1521,net_1520}),
    .q({open_n1087,net_1519})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h1000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h8800"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_728
  (
    .clk(gclk_8),
    .ce(net_1524),
    .sr(net_182),
    .a({net_1289,net_1302}),
    .b({net_1302,net_247}),
    .c({open_n1088,net_1047}),
    .d({net_963,net_948}),
    .e({net_948,net_963}),
    .mi({open_n1089,io_i2c_sda}),
    .f({net_1523,net_1524}),
    .q({open_n1090,net_1522})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h5000"),
    .INIT_LUT1("16'h0200"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_729
  (
    .clk(gclk_8),
    .ce(net_1526),
    .sr(net_182),
    .a({net_948,net_247}),
    .b({net_1182,open_n1091}),
    .c({net_1302,net_1047}),
    .d({net_1312,net_1525}),
    .mi({open_n1092,io_i2c_sda}),
    .f({net_1525,net_1526}),
    .q({open_n1093,net_1527})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h4000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("ON"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("SET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_730
  (
    .a({net_1532,net_1532}),
    .b({net_1289,net_1289}),
    .c({net_1300,net_1301}),
    .d({net_1301,net_1300}),
    .mi({open_n1094,net_1299}),
    .fx({open_n1095,net_1528})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0011"),
    .INIT_LUTG0("16'h0011"),
    .INIT_LUTF1("16'h0005"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_731
  (
    .clk(gclk_8),
    .ce(net_1530),
    .sr(net_182),
    .a({net_1529,net_1323}),
    .b({open_n1096,net_1327}),
    .c({net_1325,open_n1097}),
    .d({net_1313,net_1529}),
    .e({net_1323,open_n1098}),
    .mi({net_1315,net_1308}),
    .f({net_1531,net_1530}),
    .q({net_1529,net_1532})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h000A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_771
  (
    .clk(gclk_5),
    .sr(net_1665),
    .a({net_1559,1'b0}),
    .b({net_1589,net_1568}),
    .c({1'b0,1'b0}),
    .d({1'b0,open_n1099}),
    .e({1'b0,open_n1100}),
    .mi({net_1563,net_1567}),
    .f({net_1563,open_n1101}),
    .fx({net_1560,net_1567}),
    .q({net_1559,net_1568}),
    .fco(sig_771_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_772
  (
    .clk(gclk_5),
    .sr(net_1665),
    .a({net_1657,net_1558}),
    .b({net_1672,net_1562}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1564,net_1566}),
    .fci(sig_771_carry),
    .f({net_1565,net_1566}),
    .fx({net_1561,net_1564}),
    .q({net_1562,net_1558}),
    .fco(sig_772_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_773
  (
    .clk(gclk_5),
    .sr(net_1665),
    .a({net_1656,net_1571}),
    .b({net_1570,net_1658}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1575,net_1580}),
    .fci(sig_772_carry),
    .f({net_1573,net_1575}),
    .fx({net_1580,net_1577}),
    .q({net_1571,net_1570}),
    .fco(sig_773_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_774
  (
    .clk(gclk_5),
    .sr(net_1665),
    .a({net_1666,net_1569}),
    .b({net_1663,net_1572}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1574,net_1579}),
    .fci(sig_773_carry),
    .f({net_1578,net_1579}),
    .fx({net_1576,net_1574}),
    .q({net_1572,net_1569}),
    .fco(sig_774_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_775
  (
    .clk(gclk_5),
    .sr(net_1665),
    .a({net_1655,net_1581}),
    .b({net_1616,net_1592}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1594,net_1590}),
    .fci(sig_774_carry),
    .f({net_1591,net_1590}),
    .fx({net_1587,net_1594}),
    .q({net_1592,net_1581}),
    .fco(sig_775_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_776
  (
    .clk(gclk_5),
    .sr(net_1665),
    .a({net_1610,net_1582}),
    .b({net_1671,net_1585}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1593,net_1595}),
    .fci(sig_775_carry),
    .f({net_1586,net_1595}),
    .fx({net_1588,net_1593}),
    .q({net_1585,net_1582}),
    .fco(sig_776_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_778
  (
    .clk(gclk_5),
    .sr(net_1665),
    .a({net_1612,net_1596}),
    .b({net_1602,net_1606}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1608,net_1604}),
    .fci(sig_776_carry),
    .f({net_1599,net_1604}),
    .fx({net_1601,net_1608}),
    .q({net_1606,net_1596}),
    .fco(sig_778_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_779
  (
    .clk(gclk_5),
    .sr(net_1665),
    .a({net_1583,net_1597}),
    .b({net_1603,net_1598}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1607,net_1609}),
    .fci(sig_778_carry),
    .f({net_1600,net_1609}),
    .fx({net_1605,net_1607}),
    .q({net_1598,net_1597}),
    .fco(sig_779_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_781
  (
    .clk(gclk_5),
    .sr(net_1665),
    .a({open_n1102,net_1611}),
    .c({1'b0,1'b0}),
    .d({open_n1103,1'b0}),
    .mi({net_1587,net_1614}),
    .fci(sig_779_carry),
    .f({open_n1104,net_1614}),
    .q({net_1616,net_1611})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0100"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_777
  (
    .clk(gclk_5),
    .sr(net_1665),
    .a({open_n1105,net_1583}),
    .b({net_1347,net_1603}),
    .c({open_n1106,net_1611}),
    .d({open_n1107,net_1615}),
    .mi({net_1560,net_1600}),
    .f({open_n1108,net_1584}),
    .q({net_1589,net_1583})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_780
  (
    .clk(gclk_5),
    .sr(net_1665),
    .mi({net_1601,net_1605}),
    .q({net_1602,net_1603})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0100"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0005"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_782
  (
    .clk(gclk_5),
    .sr(net_1665),
    .a({net_1610,net_1612}),
    .b({open_n1109,net_1602}),
    .c({net_1671,net_1597}),
    .d({net_1596,net_1613}),
    .e({net_1606,net_1598}),
    .mi({net_1586,net_1599}),
    .f({net_1613,net_1615}),
    .q({net_1610,net_1612})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h5555"),
    .INIT_LUTG0("16'h5555"),
    .INIT_LUTF1("16'h5555"),
    .INIT_LUTG1("16'h5555"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("F"),
    .REG1_SD("F"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_783
  (
    .clk(gclk_0),
    .ce(net_451),
    .a({net_1618,net_1617}),
    .q({net_1618,net_1617})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h000A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_784
  (
    .clk(gclk_0),
    .sr(net_1669),
    .a({net_1620,1'b0}),
    .b({net_1667,net_1629}),
    .c({1'b0,1'b0}),
    .d({1'b0,open_n1110}),
    .e({1'b0,open_n1111}),
    .mi({net_1624,net_1628}),
    .f({net_1624,open_n1112}),
    .fx({net_1625,net_1628}),
    .q({net_1620,net_1629}),
    .fco(sig_784_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_785
  (
    .clk(gclk_0),
    .sr(net_1669),
    .a({net_1650,net_1619}),
    .b({net_1647,net_1622}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1626,net_1627}),
    .fci(sig_784_carry),
    .f({net_1621,net_1627}),
    .fx({net_1623,net_1626}),
    .q({net_1622,net_1619}),
    .fco(sig_785_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_786
  (
    .clk(gclk_0),
    .sr(net_1669),
    .a({net_1632,net_1633}),
    .b({net_1638,net_1631}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1636,net_1643}),
    .fci(sig_785_carry),
    .f({net_1637,net_1636}),
    .fx({net_1643,net_1640}),
    .q({net_1633,net_1638}),
    .fco(sig_786_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_787
  (
    .clk(gclk_0),
    .sr(net_1669),
    .a({net_1670,net_1630}),
    .b({net_1645,net_1634}),
    .c({1'b0,1'b0}),
    .d({1'b0,1'b0}),
    .e({1'b0,1'b0}),
    .mi({net_1639,net_1642}),
    .fci(sig_786_carry),
    .f({net_1641,net_1642}),
    .fx({net_1635,net_1639}),
    .q({net_1634,net_1630}),
    .fco(sig_787_carry)
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'hA55A"),
    .INIT_LUTG0("16'hC33C"),
    .INIT_LUTF1("16'hA55A"),
    .INIT_LUTG1("16'hC33C"),
    .MODE("RIPPLE"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_789
  (
    .clk(gclk_0),
    .sr(net_1669),
    .a({open_n1113,net_1644}),
    .c({1'b0,1'b0}),
    .d({open_n1114,1'b0}),
    .mi({net_1621,net_1649}),
    .fci(sig_787_carry),
    .f({open_n1115,net_1649}),
    .q({net_1650,net_1644})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0000"),
    .INIT_LUT1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_788
  (
    .clk(gclk_0),
    .sr(net_1669),
    .mi({net_1640,net_1637}),
    .q({net_1631,net_1632})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h5555"),
    .INIT_LUT1("16'h4000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("CE"),
    .SRMUX("0"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("F"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("SET"),
    .SRMODE("ASYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_790
  (
    .clk(gclk_0),
    .ce(net_1669),
    .a({net_1182,net_1646}),
    .b({net_948,open_n1116}),
    .c({net_1312,open_n1117}),
    .d({net_1302,open_n1118}),
    .f({net_1648,open_n1119}),
    .q({open_n1120,net_1646})
  );

  AL_PHY_MSLICE #
  (
    .INIT_LUT0("16'h0001"),
    .INIT_LUT1("16'h0001"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MSFXMUX("OFF"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  mslice_block_791
  (
    .clk(gclk_0),
    .sr(net_1669),
    .a({net_1645,net_1647}),
    .b({net_1644,net_1633}),
    .c({net_1634,net_1631}),
    .d({net_1670,net_1632}),
    .mi({net_1635,net_1623}),
    .f({net_1651,net_1652}),
    .q({net_1645,net_1647})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0101"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'hDF00"),
    .INIT_LUTG1("16'hDF00"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_796
  (
    .clk(gclk_5),
    .sr(net_1665),
    .a({net_1658,net_1656}),
    .b({net_1660,net_1569}),
    .c({net_1571,net_1572}),
    .d({net_1659,open_n1121}),
    .e({open_n1122,net_1570}),
    .mi({net_1577,net_1573}),
    .f({net_1661,net_1659}),
    .q({net_1658,net_1656})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0077"),
    .INIT_LUTG0("16'h0055"),
    .INIT_LUTF1("16'h0101"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_797
  (
    .clk(gclk_5),
    .sr(net_1665),
    .a({net_1655,net_1657}),
    .b({net_1616,net_1562}),
    .c({net_1582,open_n1123}),
    .d({open_n1124,net_1672}),
    .e({net_1585,net_1558}),
    .mi({net_1591,net_1565}),
    .f({net_1662,net_1660}),
    .q({net_1655,net_1657})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h7555"),
    .INIT_LUTG0("16'h7555"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h000C"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_798
  (
    .clk(gclk_5),
    .sr(net_1665),
    .a({open_n1125,net_1664}),
    .b({net_1584,net_1661}),
    .c({net_1581,net_1666}),
    .d({net_1592,net_1663}),
    .e({net_1662,open_n1126}),
    .mi({net_1576,net_1578}),
    .f({net_1664,net_1665}),
    .q({net_1663,net_1666})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h7FFF"),
    .INIT_LUTF1("16'hDDFF"),
    .INIT_LUTG1("16'hFFFF"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_799
  (
    .clk(gclk_0),
    .sr(net_1669),
    .a({net_1668,net_1667}),
    .b({net_1630,net_1622}),
    .c({open_n1127,net_1650}),
    .d({net_1651,net_1619}),
    .e({net_1638,net_1652}),
    .mi({net_1641,net_1625}),
    .f({net_1669,net_1668}),
    .q({net_1670,net_1667})
  );

  AL_PHY_LSLICE #
  (
    .INIT_LUTF0("16'h0000"),
    .INIT_LUTG0("16'h0000"),
    .INIT_LUTF1("16'h0000"),
    .INIT_LUTG1("16'h0000"),
    .MODE("LOGIC"),
    .GSR("ENABLE"),
    .CEMUX("1"),
    .SRMUX("SR"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .DEMUX0("D"),
    .DEMUX1("D"),
    .CMIMUX0("C"),
    .CMIMUX1("C"),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .LSFXMUX0("FUNC5"),
    .LSFXMUX1("FUNC5"),
    .REG0_SD("MI"),
    .REG1_SD("MI"),
    .REG0_REGSET("RESET"),
    .REG1_REGSET("RESET"),
    .SRMODE("SYNC"),
    .TESTMODE("OFF")
  )
  lslice_block_800
  (
    .clk(gclk_5),
    .sr(net_1665),
    .mi({net_1588,net_1561}),
    .q({net_1671,net_1672})
  );

  AL_PHY_BRAM #
  (
    //.RID("0x0004"),
    //.WID("0x0004"),
    .MODE("DP8K"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("READBEFOREWRITE"),
    .GSR("ENABLE"),
    .RESETMODE("ASYNC"),
    .ASYNC_RESET_RELEASE("SYNC"),
    .CEAMUX("0"),
    .CEBMUX("0"),
    .OCEAMUX("SIG"),
    .OCEBMUX("SIG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .CLKAMUX("SIG"),
    .CLKBMUX("SIG"),
    .WEAMUX("0"),
    .WEBMUX("SIG"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1")
  )
  emb_block_61
  (
    .dia({open_n1128,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
    .doa({open_n1129,net_28,net_25,net_26,net_27,net_24,net_21,net_23,net_22}),
    .addra({net_76,net_74,net_77,net_70,net_72,net_71,net_73,net_67,net_69,net_68,open_n1130,open_n1131,open_n1132}),
    .csa({1'b0,1'b0,1'b0}),
    .clka(gclk_7),
    .dib({open_n1133,io_mcu_d[7],io_mcu_d[6],io_mcu_d[5],io_mcu_d[4],io_mcu_d[3],io_mcu_d[2],io_mcu_d[1],io_mcu_d[0]}),
    .addrb({net_126,net_128,net_130,net_119,net_118,net_117,net_120,net_111,net_110,net_112,open_n1134,open_n1135,open_n1136}),
    .csb({1'b0,1'b0,1'b0}),
    .web(net_512),
    .clkb(gclk_9)
  );

  AL_PHY_BRAM #
  (
    //.RID("0x000E"),
    //.WID("0x000E"),
    .MODE("DP8K"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .WRITEMODE_A("WRITETHROUGH"),
    .WRITEMODE_B("READBEFOREWRITE"),
    .GSR("ENABLE"),
    .RESETMODE("SYNC"),
    .ASYNC_RESET_RELEASE("SYNC"),
    .CEAMUX("SIG"),
    .CEBMUX("0"),
    .OCEAMUX("SIG"),
    .OCEBMUX("SIG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .CLKAMUX("SIG"),
    .CLKBMUX("SIG"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("1")
  )
  emb_block_69
  (
    .dia({net_1007,net_819,net_933,net_1237,net_1046,net_799,net_1250,net_1011,net_1139}),
    .addra({net_872,net_988,net_1211,net_986,net_992,net_1096,net_1006,net_1103,net_1511,net_1219,open_n1137,open_n1138,open_n1139}),
    .csa({1'b0,net_1133,net_1218}),
    .cea(net_1496),
    .clka(gclk_4),
    .dob({net_33,net_37,net_35,net_36,net_34,net_30,net_29,net_31,net_32}),
    .addrb({net_1294,net_1298,net_1154,net_1147,net_1031,net_921,net_924,net_1146,net_1290,net_1512,open_n1140,open_n1141,open_n1142}),
    .csb({1'b0,net_193,net_1050}),
    .clkb(gclk_3)
  );

  AL_PHY_BRAM #
  (
    //.RID("0x0011"),
    //.WID("0x0011"),
    .MODE("DP8K"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .WRITEMODE_A("WRITETHROUGH"),
    .WRITEMODE_B("READBEFOREWRITE"),
    .GSR("ENABLE"),
    .RESETMODE("SYNC"),
    .ASYNC_RESET_RELEASE("SYNC"),
    .CEAMUX("SIG"),
    .CEBMUX("0"),
    .OCEAMUX("SIG"),
    .OCEBMUX("SIG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .CLKAMUX("SIG"),
    .CLKBMUX("SIG"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("1")
  )
  emb_block_70
  (
    .dia({net_1007,net_819,net_933,net_1237,net_1046,net_799,net_1250,net_1011,net_1139}),
    .addra({net_872,net_988,net_1211,net_986,net_992,net_1096,net_1006,net_1103,net_1511,net_1219,open_n1143,open_n1144,open_n1145}),
    .csa({1'b0,net_1133,net_1218}),
    .cea(net_1496),
    .clka(gclk_4),
    .dob({net_43,net_46,net_42,net_45,net_44,net_41,net_38,net_39,net_40}),
    .addrb({net_1294,net_1298,net_1154,net_1147,net_1031,net_921,net_924,net_1146,net_1290,net_1512,open_n1146,open_n1147,open_n1148}),
    .csb({1'b0,net_193,net_1050}),
    .clkb(gclk_3)
  );

  AL_PHY_BRAM #
  (
    //.RID("0x0005"),
    //.WID("0x0005"),
    .MODE("DP8K"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .WRITEMODE_A("WRITETHROUGH"),
    .WRITEMODE_B("READBEFOREWRITE"),
    .GSR("ENABLE"),
    .RESETMODE("SYNC"),
    .ASYNC_RESET_RELEASE("SYNC"),
    .CEAMUX("SIG"),
    .CEBMUX("0"),
    .OCEAMUX("SIG"),
    .OCEBMUX("SIG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .CLKAMUX("SIG"),
    .CLKBMUX("SIG"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("1")
  )
  emb_block_71
  (
    .dia({net_1007,net_819,net_933,net_1237,net_1046,net_799,net_1250,net_1011,net_1139}),
    .addra({net_872,net_988,net_1211,net_986,net_992,net_1096,net_1006,net_1103,net_1511,net_1219,open_n1149,open_n1150,open_n1151}),
    .csa({1'b0,net_1133,net_1218}),
    .cea(net_1496),
    .clka(gclk_4),
    .dob({net_52,net_53,net_51,net_55,net_54,net_47,net_48,net_49,net_50}),
    .addrb({net_1294,net_1298,net_1154,net_1147,net_1031,net_921,net_924,net_1146,net_1290,net_1512,open_n1152,open_n1153,open_n1154}),
    .csb({1'b0,net_193,net_1050}),
    .clkb(gclk_3)
  );

  AL_PHY_BRAM #
  (
    //.RID("0x000B"),
    //.WID("0x000B"),
    .MODE("DP8K"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .WRITEMODE_A("WRITETHROUGH"),
    .WRITEMODE_B("READBEFOREWRITE"),
    .GSR("ENABLE"),
    .RESETMODE("SYNC"),
    .ASYNC_RESET_RELEASE("SYNC"),
    .CEAMUX("SIG"),
    .CEBMUX("0"),
    .OCEAMUX("SIG"),
    .OCEBMUX("SIG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .CLKAMUX("SIG"),
    .CLKBMUX("SIG"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("1")
  )
  emb_block_88
  (
    .dia({net_1007,net_819,net_933,net_1237,net_1046,net_799,net_1250,net_1011,net_1139}),
    .addra({net_872,net_988,net_1211,net_986,net_992,net_1096,net_1006,net_1103,net_1511,net_1219,open_n1155,open_n1156,open_n1157}),
    .csa({1'b0,net_1133,net_1218}),
    .cea(net_1496),
    .clka(gclk_4),
    .dob({net_58,net_64,net_61,net_63,net_62,net_56,net_57,net_60,net_59}),
    .addrb({net_1294,net_1298,net_1154,net_1147,net_1031,net_921,net_924,net_1146,net_1290,net_1512,open_n1158,open_n1159,open_n1160}),
    .csb({1'b0,net_193,net_1050}),
    .clkb(gclk_3)
  );

  AL_PHY_BRAM #
  (
    //.RID("0x0007"),
    //.WID("0x0007"),
    .MODE("DP8K"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .WRITEMODE_A("WRITETHROUGH"),
    .WRITEMODE_B("READBEFOREWRITE"),
    .GSR("ENABLE"),
    .RESETMODE("SYNC"),
    .ASYNC_RESET_RELEASE("SYNC"),
    .CEAMUX("SIG"),
    .CEBMUX("0"),
    .OCEAMUX("SIG"),
    .OCEBMUX("SIG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .CLKAMUX("SIG"),
    .CLKBMUX("SIG"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("1")
  )
  emb_block_390
  (
    .dia({net_1254,net_1012,net_1246,net_1489,net_1504,net_1236,net_1487,net_1340,net_1248}),
    .addra({net_872,net_988,net_1211,net_986,net_992,net_1096,net_1006,net_1103,net_1511,net_1219,open_n1161,open_n1162,open_n1163}),
    .csa({1'b0,net_1133,net_1218}),
    .cea(net_1496),
    .clka(gclk_4),
    .dob({net_690,net_697,net_696,net_698,net_695,net_693,net_694,net_691,net_692}),
    .addrb({net_1294,net_1298,net_1154,net_1147,net_1031,net_921,net_924,net_1146,net_1290,net_1512,open_n1164,open_n1165,open_n1166}),
    .csb({1'b0,net_193,net_1050}),
    .clkb(gclk_3)
  );

  AL_PHY_BRAM #
  (
    //.RID("0x000D"),
    //.WID("0x000D"),
    .MODE("DP8K"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .WRITEMODE_A("WRITETHROUGH"),
    .WRITEMODE_B("READBEFOREWRITE"),
    .GSR("ENABLE"),
    .RESETMODE("SYNC"),
    .ASYNC_RESET_RELEASE("SYNC"),
    .CEAMUX("SIG"),
    .CEBMUX("0"),
    .OCEAMUX("SIG"),
    .OCEBMUX("SIG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .CLKAMUX("SIG"),
    .CLKBMUX("SIG"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("1")
  )
  emb_block_398
  (
    .dia({net_1254,net_1012,net_1246,net_1489,net_1504,net_1236,net_1487,net_1340,net_1248}),
    .addra({net_872,net_988,net_1211,net_986,net_992,net_1096,net_1006,net_1103,net_1511,net_1219,open_n1167,open_n1168,open_n1169}),
    .csa({1'b0,net_1133,net_1218}),
    .cea(net_1496),
    .clka(gclk_4),
    .dob({net_702,net_705,net_706,net_704,net_707,net_703,net_699,net_701,net_700}),
    .addrb({net_1294,net_1298,net_1154,net_1147,net_1031,net_921,net_924,net_1146,net_1290,net_1512,open_n1170,open_n1171,open_n1172}),
    .csb({1'b0,net_193,net_1050}),
    .clkb(gclk_3)
  );

  AL_PHY_BRAM #
  (
    //.RID("0x000F"),
    //.WID("0x000F"),
    .MODE("DP8K"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .WRITEMODE_A("WRITETHROUGH"),
    .WRITEMODE_B("READBEFOREWRITE"),
    .GSR("ENABLE"),
    .RESETMODE("SYNC"),
    .ASYNC_RESET_RELEASE("SYNC"),
    .CEAMUX("SIG"),
    .CEBMUX("0"),
    .OCEAMUX("SIG"),
    .OCEBMUX("SIG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .CLKAMUX("SIG"),
    .CLKBMUX("SIG"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("1")
  )
  emb_block_399
  (
    .dia({net_806,net_1257,net_1104,net_938,net_818,net_1051,net_1134,net_1517,net_944}),
    .addra({net_872,net_988,net_1211,net_986,net_992,net_1096,net_1006,net_1103,net_1511,net_1219,open_n1173,open_n1174,open_n1175}),
    .csa({1'b0,net_1133,net_1218}),
    .cea(net_1496),
    .clka(gclk_4),
    .dob({net_712,net_714,net_715,net_716,net_713,net_711,net_708,net_710,net_709}),
    .addrb({net_1294,net_1298,net_1154,net_1147,net_1031,net_921,net_924,net_1146,net_1290,net_1512,open_n1176,open_n1177,open_n1178}),
    .csb({1'b0,net_193,net_1050}),
    .clkb(gclk_3)
  );

  AL_PHY_BRAM #
  (
    //.RID("0x0012"),
    //.WID("0x0012"),
    .MODE("DP8K"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .WRITEMODE_A("WRITETHROUGH"),
    .WRITEMODE_B("READBEFOREWRITE"),
    .GSR("ENABLE"),
    .RESETMODE("SYNC"),
    .ASYNC_RESET_RELEASE("SYNC"),
    .CEAMUX("SIG"),
    .CEBMUX("0"),
    .OCEAMUX("SIG"),
    .OCEBMUX("SIG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .CLKAMUX("SIG"),
    .CLKBMUX("SIG"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("1")
  )
  emb_block_400
  (
    .dia({net_806,net_1257,net_1104,net_938,net_818,net_1051,net_1134,net_1517,net_944}),
    .addra({net_872,net_988,net_1211,net_986,net_992,net_1096,net_1006,net_1103,net_1511,net_1219,open_n1179,open_n1180,open_n1181}),
    .csa({1'b0,net_1133,net_1218}),
    .cea(net_1496),
    .clka(gclk_4),
    .dob({net_722,net_725,net_721,net_723,net_724,net_717,net_720,net_718,net_719}),
    .addrb({net_1294,net_1298,net_1154,net_1147,net_1031,net_921,net_924,net_1146,net_1290,net_1512,open_n1182,open_n1183,open_n1184}),
    .csb({1'b0,net_193,net_1050}),
    .clkb(gclk_3)
  );

  AL_PHY_BRAM #
  (
    //.RID("0x000C"),
    //.WID("0x000C"),
    .MODE("DP8K"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .WRITEMODE_A("WRITETHROUGH"),
    .WRITEMODE_B("READBEFOREWRITE"),
    .GSR("ENABLE"),
    .RESETMODE("SYNC"),
    .ASYNC_RESET_RELEASE("SYNC"),
    .CEAMUX("SIG"),
    .CEBMUX("0"),
    .OCEAMUX("SIG"),
    .OCEBMUX("SIG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .CLKAMUX("SIG"),
    .CLKBMUX("SIG"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("1")
  )
  emb_block_401
  (
    .dia({net_806,net_1257,net_1104,net_938,net_818,net_1051,net_1134,net_1517,net_944}),
    .addra({net_872,net_988,net_1211,net_986,net_992,net_1096,net_1006,net_1103,net_1511,net_1219,open_n1185,open_n1186,open_n1187}),
    .csa({1'b0,net_1133,net_1218}),
    .cea(net_1496),
    .clka(gclk_4),
    .dob({net_728,net_732,net_733,net_734,net_731,net_730,net_729,net_727,net_726}),
    .addrb({net_1294,net_1298,net_1154,net_1147,net_1031,net_921,net_924,net_1146,net_1290,net_1512,open_n1188,open_n1189,open_n1190}),
    .csb({1'b0,net_193,net_1050}),
    .clkb(gclk_3)
  );

  AL_PHY_BRAM #
  (
    //.RID("0x0006"),
    //.WID("0x0006"),
    .MODE("DP8K"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .WRITEMODE_A("WRITETHROUGH"),
    .WRITEMODE_B("READBEFOREWRITE"),
    .GSR("ENABLE"),
    .RESETMODE("SYNC"),
    .ASYNC_RESET_RELEASE("SYNC"),
    .CEAMUX("SIG"),
    .CEBMUX("0"),
    .OCEAMUX("SIG"),
    .OCEBMUX("SIG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .CLKAMUX("SIG"),
    .CLKBMUX("SIG"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("1")
  )
  emb_block_406
  (
    .dia({net_806,net_1257,net_1104,net_938,net_818,net_1051,net_1134,net_1517,net_944}),
    .addra({net_872,net_988,net_1211,net_986,net_992,net_1096,net_1006,net_1103,net_1511,net_1219,open_n1191,open_n1192,open_n1193}),
    .csa({1'b0,net_1133,net_1218}),
    .cea(net_1496),
    .clka(gclk_4),
    .dob({net_738,net_741,net_743,net_740,net_742,net_739,net_737,net_736,net_735}),
    .addrb({net_1294,net_1298,net_1154,net_1147,net_1031,net_921,net_924,net_1146,net_1290,net_1512,open_n1194,open_n1195,open_n1196}),
    .csb({1'b0,net_193,net_1050}),
    .clkb(gclk_3)
  );

  AL_PHY_BRAM #
  (
    //.RID("0x0010"),
    //.WID("0x0010"),
    .MODE("DP8K"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .WRITEMODE_A("WRITETHROUGH"),
    .WRITEMODE_B("READBEFOREWRITE"),
    .GSR("ENABLE"),
    .RESETMODE("SYNC"),
    .ASYNC_RESET_RELEASE("SYNC"),
    .CEAMUX("SIG"),
    .CEBMUX("0"),
    .OCEAMUX("SIG"),
    .OCEBMUX("SIG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .CLKAMUX("SIG"),
    .CLKBMUX("SIG"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("1")
  )
  emb_block_732
  (
    .dia({net_1254,net_1012,net_1246,net_1489,net_1504,net_1236,net_1487,net_1340,net_1248}),
    .addra({net_872,net_988,net_1211,net_986,net_992,net_1096,net_1006,net_1103,net_1511,net_1219,open_n1197,open_n1198,open_n1199}),
    .csa({1'b0,net_1133,net_1218}),
    .cea(net_1496),
    .clka(gclk_4),
    .dob({net_1534,net_1540,net_1542,net_1539,net_1541,net_1537,net_1538,net_1535,net_1536}),
    .addrb({net_1294,net_1298,net_1154,net_1147,net_1031,net_921,net_924,net_1146,net_1290,net_1512,open_n1200,open_n1201,open_n1202}),
    .csb({1'b0,net_193,net_1050}),
    .clkb(gclk_3)
  );

  AL_PHY_BRAM #
  (
    //.RID("0x0013"),
    //.WID("0x0013"),
    .MODE("DP8K"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .WRITEMODE_A("WRITETHROUGH"),
    .WRITEMODE_B("READBEFOREWRITE"),
    .GSR("ENABLE"),
    .RESETMODE("SYNC"),
    .ASYNC_RESET_RELEASE("SYNC"),
    .CEAMUX("SIG"),
    .CEBMUX("0"),
    .OCEAMUX("SIG"),
    .OCEBMUX("SIG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .CLKAMUX("SIG"),
    .CLKBMUX("SIG"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("1")
  )
  emb_block_738
  (
    .dia({net_1254,net_1012,net_1246,net_1489,net_1504,net_1236,net_1487,net_1340,net_1248}),
    .addra({net_872,net_988,net_1211,net_986,net_992,net_1096,net_1006,net_1103,net_1511,net_1219,open_n1203,open_n1204,open_n1205}),
    .csa({1'b0,net_1133,net_1218}),
    .cea(net_1496),
    .clka(gclk_4),
    .dob({net_1544,net_1549,net_1550,net_1548,net_1551,net_1546,net_1545,net_1543,net_1547}),
    .addrb({net_1294,net_1298,net_1154,net_1147,net_1031,net_921,net_924,net_1146,net_1290,net_1512,open_n1206,open_n1207,open_n1208}),
    .csb({1'b0,net_193,net_1050}),
    .clkb(gclk_3)
  );

  AL_PHY_BRAM #
  (
    //.RID("0x000A"),
    //.WID("0x000A"),
    .MODE("DP8K"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .WRITEMODE_A("WRITETHROUGH"),
    .WRITEMODE_B("READBEFOREWRITE"),
    .GSR("ENABLE"),
    .RESETMODE("SYNC"),
    .ASYNC_RESET_RELEASE("SYNC"),
    .CEAMUX("SIG"),
    .CEBMUX("0"),
    .OCEAMUX("SIG"),
    .OCEBMUX("SIG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .CLKAMUX("SIG"),
    .CLKBMUX("SIG"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1")
  )
  emb_block_739
  (
    .dia({open_n1209,open_n1210,open_n1211,open_n1212,open_n1213,open_n1214,net_1488,open_n1215,open_n1216}),
    .addra({net_1133,net_1218,net_872,net_988,net_1211,net_986,net_992,net_1096,net_1006,net_1103,net_1511,net_1219,open_n1217}),
    .csa({1'b0,1'b0,1'b0}),
    .cea(net_1496),
    .clka(gclk_4),
    .dob({open_n1218,open_n1219,open_n1220,open_n1221,open_n1222,open_n1223,open_n1224,open_n1225,net_1552}),
    .addrb({net_193,net_1050,net_1294,net_1298,net_1154,net_1147,net_1031,net_921,net_924,net_1146,net_1290,net_1512,open_n1226}),
    .csb({1'b0,1'b0,1'b0}),
    .clkb(gclk_3)
  );

  AL_PHY_BRAM #
  (
    //.RID("0x0008"),
    //.WID("0x0008"),
    .MODE("DP8K"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .WRITEMODE_A("WRITETHROUGH"),
    .WRITEMODE_B("READBEFOREWRITE"),
    .GSR("ENABLE"),
    .RESETMODE("SYNC"),
    .ASYNC_RESET_RELEASE("SYNC"),
    .CEAMUX("SIG"),
    .CEBMUX("0"),
    .OCEAMUX("SIG"),
    .OCEBMUX("SIG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .CLKAMUX("SIG"),
    .CLKBMUX("SIG"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1")
  )
  emb_block_740
  (
    .dia({open_n1227,open_n1228,open_n1229,net_1486,open_n1230,open_n1231,net_1346,open_n1232,open_n1233}),
    .addra({net_1133,net_1218,net_872,net_988,net_1211,net_986,net_992,net_1096,net_1006,net_1103,net_1511,net_1219,open_n1234}),
    .csa({1'b0,1'b0,1'b0}),
    .cea(net_1496),
    .clka(gclk_4),
    .dob({open_n1235,open_n1236,open_n1237,open_n1238,open_n1239,open_n1240,open_n1241,net_1553,net_1554}),
    .addrb({net_193,net_1050,net_1294,net_1298,net_1154,net_1147,net_1031,net_921,net_924,net_1146,net_1290,net_1512,open_n1242}),
    .csb({1'b0,1'b0,1'b0}),
    .clkb(gclk_3)
  );

  AL_PHY_BRAM #
  (
    //.RID("0x0009"),
    //.WID("0x0009"),
    .MODE("DP8K"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .WRITEMODE_A("WRITETHROUGH"),
    .WRITEMODE_B("READBEFOREWRITE"),
    .GSR("ENABLE"),
    .RESETMODE("SYNC"),
    .ASYNC_RESET_RELEASE("SYNC"),
    .CEAMUX("SIG"),
    .CEBMUX("0"),
    .OCEAMUX("SIG"),
    .OCEBMUX("SIG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .CLKAMUX("SIG"),
    .CLKBMUX("SIG"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1")
  )
  emb_block_757
  (
    .dia({open_n1243,open_n1244,open_n1245,net_1506,open_n1246,open_n1247,net_1243,open_n1248,open_n1249}),
    .addra({net_1133,net_1218,net_872,net_988,net_1211,net_986,net_992,net_1096,net_1006,net_1103,net_1511,net_1219,open_n1250}),
    .csa({1'b0,1'b0,1'b0}),
    .cea(net_1496),
    .clka(gclk_4),
    .dob({open_n1251,open_n1252,open_n1253,open_n1254,open_n1255,open_n1256,open_n1257,net_1555,net_1556}),
    .addrb({net_193,net_1050,net_1294,net_1298,net_1154,net_1147,net_1031,net_921,net_924,net_1146,net_1290,net_1512,open_n1258}),
    .csb({1'b0,1'b0,1'b0}),
    .clkb(gclk_3)
  );

  AL_PHY_PLL #
  (
    .FIN("50.000"),
    .FEEDBK_MODE("NOCOMP"),
    .FEEDBK_PATH("VCO_PHASE_0"),
    .STDBY_ENABLE("DISABLE"),
    .PLLRST_ENA("ENABLE"),
    .SYNC_ENABLE("DISABLE"),
    .DERIVE_PLL_CLOCKS("DISABLE"),
    .GEN_BASIC_CLOCK("DISABLE"),
    .GMC_GAIN("4"),
    .ICP_CURRENT(11),
    .KVCO("4"),
    .LPF_CAPACITOR("1"),
    .LPF_RESISTOR(4),
    .REFCLK_DIV(1),
    .FBCLK_DIV(20),
    .CLKC0_ENABLE("ENABLE"),
    .CLKC0_DIV(5),
    .CLKC0_CPHASE(4),
    .CLKC0_FPHASE("0")
  )
  pll_inst
  (
    .refclk(i_xtal),
    .pllreset(1'b0),
    .stdby(1'b0),
    .ext_lock(open),
    .load_reg(1'b0),
    .scanclk(1'b0),
    .phaseupdown(1'b0),
    .phasestep(1'b0),
    .phcntsel(3'b000),
    .phasedone(open),
    .fbclk(1'b0),
    .clkc({open, open, open, open, clock_200MHz})
  );

endmodule

